module vscale_core ( clk, ext_interrupts, imem_haddr, imem_hwrite, imem_hsize, 
        imem_hburst, imem_hmastlock, imem_hprot, imem_htrans, imem_hwdata, 
        imem_hrdata, imem_hready, imem_hresp, dmem_haddr, dmem_hwrite, 
        dmem_hsize, dmem_hburst, dmem_hmastlock, dmem_hprot, dmem_htrans, 
        dmem_hwdata, dmem_hrdata, dmem_hready, dmem_hresp, htif_reset, htif_id, 
        htif_pcr_req_valid, htif_pcr_req_ready, htif_pcr_req_rw, 
        htif_pcr_req_addr, htif_pcr_req_data, htif_pcr_resp_valid, 
        htif_pcr_resp_ready, htif_pcr_resp_data, htif_ipi_req_ready, 
        htif_ipi_req_valid, htif_ipi_req_data, htif_ipi_resp_ready, 
        htif_ipi_resp_valid, htif_ipi_resp_data, htif_debug_stats_pcr );
  input [23:0] ext_interrupts;
  output [31:0] imem_haddr;
  output [2:0] imem_hsize;
  output [2:0] imem_hburst;
  output [3:0] imem_hprot;
  output [1:0] imem_htrans;
  output [31:0] imem_hwdata;
  input [31:0] imem_hrdata;
  input imem_hresp;
  output [31:0] dmem_haddr;
  output [2:0] dmem_hsize;
  output [2:0] dmem_hburst;
  output [3:0] dmem_hprot;
  output [1:0] dmem_htrans;
  output [31:0] dmem_hwdata;
  input [31:0] dmem_hrdata;
  input dmem_hresp;
  input [11:0] htif_pcr_req_addr;
  input [63:0] htif_pcr_req_data;
  output [63:0] htif_pcr_resp_data;
  input clk, imem_hready, dmem_hready, htif_reset, htif_id, htif_pcr_req_valid,
         htif_pcr_req_rw, htif_pcr_resp_ready, htif_ipi_req_ready,
         htif_ipi_resp_valid, htif_ipi_resp_data, pipeline_csr_system_wen, pipeline_csr_N2405, pipeline_csr_N2407;
  output imem_hwrite, imem_hmastlock, dmem_hwrite, dmem_hmastlock,
         htif_pcr_req_ready, htif_pcr_resp_valid, htif_ipi_req_valid,
         htif_ipi_req_data, htif_ipi_resp_ready, htif_debug_stats_pcr;
  wire   n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, pipeline_store_data_WB_31_, pipeline_imm_31_,
         pipeline_PC_IF_8_, pipeline_wb_src_sel_WB_0_, pipeline_dmem_type_2_,
         pipeline_ctrl_dmem_en_WB, pipeline_ctrl_wr_reg_unkilled_WB,
         pipeline_ctrl_had_ex_WB, pipeline_ctrl_N82, pipeline_ctrl_N81,
         pipeline_ctrl_prev_killed_DX, pipeline_ctrl_had_ex_DX,
         pipeline_ctrl_N66, pipeline_ctrl_replay_IF, pipeline_regfile_N21,
         pipeline_regfile_N20, pipeline_regfile_N19, pipeline_regfile_N18,
         pipeline_regfile_N17, pipeline_regfile_N16, pipeline_regfile_N15,
         pipeline_regfile_N14, pipeline_regfile_N13, pipeline_regfile_N12,
         pipeline_alu_N320, pipeline_alu_N319, pipeline_alu_N316,
         pipeline_alu_N284, pipeline_alu_N283, pipeline_alu_N282,
         pipeline_alu_N281, pipeline_alu_N280, pipeline_alu_N279,
         pipeline_alu_N278, pipeline_alu_N277, pipeline_alu_N276,
         pipeline_alu_N275, pipeline_alu_N274, pipeline_alu_N273,
         pipeline_alu_N272, pipeline_alu_N271, pipeline_alu_N270,
         pipeline_alu_N269, pipeline_alu_N268, pipeline_alu_N267,
         pipeline_alu_N266, pipeline_alu_N265, pipeline_alu_N264,
         pipeline_alu_N263, pipeline_alu_N262, pipeline_alu_N261,
         pipeline_alu_N260, pipeline_alu_N259, pipeline_alu_N258,
         pipeline_alu_N257, pipeline_alu_N256, pipeline_alu_N255,
         pipeline_alu_N254, pipeline_alu_N253, pipeline_alu_N252,
         pipeline_alu_N251, pipeline_alu_N90, pipeline_alu_N89,
         pipeline_alu_N88, pipeline_alu_N87, pipeline_alu_N86,
         pipeline_alu_N85, pipeline_alu_N84, pipeline_alu_N83,
         pipeline_alu_N82, pipeline_alu_N81, pipeline_alu_N80,
         pipeline_alu_N79, pipeline_alu_N78, pipeline_alu_N77,
         pipeline_alu_N76, pipeline_alu_N75, pipeline_alu_N74,
         pipeline_alu_N73, pipeline_alu_N72, pipeline_alu_N71,
         pipeline_alu_N70, pipeline_alu_N69, pipeline_alu_N68,
         pipeline_alu_N67, pipeline_alu_N66, pipeline_alu_N65,
         pipeline_alu_N64, pipeline_alu_N63, pipeline_alu_N62,
         pipeline_alu_N61, pipeline_alu_N60, pipeline_alu_N59,
         pipeline_md_N346, pipeline_md_N345, pipeline_md_N344,
         pipeline_md_N343, pipeline_md_N342, pipeline_md_N341,
         pipeline_md_N340, pipeline_md_N339, pipeline_md_N338,
         pipeline_md_N337, pipeline_md_N336, pipeline_md_N335,
         pipeline_md_N334, pipeline_md_N333, pipeline_md_N332,
         pipeline_md_N331, pipeline_md_N330, pipeline_md_N329,
         pipeline_md_N328, pipeline_md_N327, pipeline_md_N326,
         pipeline_md_N325, pipeline_md_N324, pipeline_md_N323,
         pipeline_md_N322, pipeline_md_N321, pipeline_md_N320,
         pipeline_md_N319, pipeline_md_N318, pipeline_md_N317,
         pipeline_md_N316, pipeline_md_N315, pipeline_md_N314,
         pipeline_md_N313, pipeline_md_N312, pipeline_md_N311,
         pipeline_md_N310, pipeline_md_N309, pipeline_md_N308,
         pipeline_md_N307, pipeline_md_N306, pipeline_md_N305,
         pipeline_md_N304, pipeline_md_N303, pipeline_md_N302,
         pipeline_md_N301, pipeline_md_N300, pipeline_md_N299,
         pipeline_md_N298, pipeline_md_N297, pipeline_md_N296,
         pipeline_md_N295, pipeline_md_N294, pipeline_md_N293,
         pipeline_md_N292, pipeline_md_N291, pipeline_md_N290,
         pipeline_md_N289, pipeline_md_N288, pipeline_md_N287,
         pipeline_md_N286, pipeline_md_N285, pipeline_md_N284,
         pipeline_md_N283, pipeline_md_N282, pipeline_md_N281,
         pipeline_md_N280, pipeline_md_N279, pipeline_md_N278,
         pipeline_md_N277, pipeline_md_N276, pipeline_md_N275,
         pipeline_md_N274, pipeline_md_N273, pipeline_md_N272,
         pipeline_md_N271, pipeline_md_N270, pipeline_md_N269,
         pipeline_md_N268, pipeline_md_N267, pipeline_md_N266,
         pipeline_md_N265, pipeline_md_N264, pipeline_md_N263,
         pipeline_md_N262, pipeline_md_N261, pipeline_md_N260,
         pipeline_md_N259, pipeline_md_N258, pipeline_md_N257,
         pipeline_md_N256, pipeline_md_N255, pipeline_md_N254,
         pipeline_md_N253, pipeline_md_N252, pipeline_md_N251,
         pipeline_md_N249, pipeline_md_N248, pipeline_md_N247,
         pipeline_md_N246, pipeline_md_N245, pipeline_md_N244,
         pipeline_md_N243, pipeline_md_N242, pipeline_md_N241,
         pipeline_md_N240, pipeline_md_N239, pipeline_md_N238,
         pipeline_md_N237, pipeline_md_N236, pipeline_md_N235,
         pipeline_md_N234, pipeline_md_N233, pipeline_md_N232,
         pipeline_md_N231, pipeline_md_N230, pipeline_md_N229,
         pipeline_md_N228, pipeline_md_N227, pipeline_md_N226,
         pipeline_md_N225, pipeline_md_N224, pipeline_md_N223,
         pipeline_md_N222, pipeline_md_N221, pipeline_md_N220,
         pipeline_md_N219, pipeline_md_N218, pipeline_md_N217,
         pipeline_md_N216, pipeline_md_N215, pipeline_md_N214,
         pipeline_md_N213, pipeline_md_N212, pipeline_md_N211,
         pipeline_md_N210, pipeline_md_N209, pipeline_md_N208,
         pipeline_md_N207, pipeline_md_N206, pipeline_md_N205,
         pipeline_md_N204, pipeline_md_N203, pipeline_md_N202,
         pipeline_md_N201, pipeline_md_N200, pipeline_md_N199,
         pipeline_md_N198, pipeline_md_N197, pipeline_md_N196,
         pipeline_md_N195, pipeline_md_N194, pipeline_md_N193,
         pipeline_md_N192, pipeline_md_N191, pipeline_md_N190,
         pipeline_md_N189, pipeline_md_N188, pipeline_md_N187,
         pipeline_md_N186, pipeline_md_N185, pipeline_md_N183,
         pipeline_md_N182, pipeline_md_N181, pipeline_md_op_0_,
         pipeline_md_N162, pipeline_md_N161, pipeline_md_N159,
         pipeline_md_N158, pipeline_md_N157, pipeline_md_N156,
         pipeline_md_N155, pipeline_md_N154, pipeline_md_N153,
         pipeline_md_N152, pipeline_md_N151, pipeline_md_N150,
         pipeline_md_N149, pipeline_md_N148, pipeline_md_N147,
         pipeline_md_N146, pipeline_md_N145, pipeline_md_N144,
         pipeline_md_N143, pipeline_md_N142, pipeline_md_N141,
         pipeline_md_N140, pipeline_md_N139, pipeline_md_N138,
         pipeline_md_N137, pipeline_md_N136, pipeline_md_N135,
         pipeline_md_N134, pipeline_md_N133, pipeline_md_N132,
         pipeline_md_N131, pipeline_md_N130, pipeline_md_N129,
         pipeline_md_N128, pipeline_md_N127, pipeline_md_N126,
         pipeline_md_N125, pipeline_md_N124, pipeline_md_N123,
         pipeline_md_N122, pipeline_md_N121, pipeline_md_N120,
         pipeline_md_N119, pipeline_md_N118, pipeline_md_N117,
         pipeline_md_N116, pipeline_md_N115, pipeline_md_N114,
         pipeline_md_N113, pipeline_md_N112, pipeline_md_N111,
         pipeline_md_N110, pipeline_md_N109, pipeline_md_N108,
         pipeline_md_N107, pipeline_md_N106, pipeline_md_N105,
         pipeline_md_N104, pipeline_md_N103, pipeline_md_N102,
         pipeline_md_N101, pipeline_md_N100, pipeline_md_N99, pipeline_md_N98,
         pipeline_md_N97, pipeline_md_N96, pipeline_md_a_geq, pipeline_md_N94,
         pipeline_md_N93, pipeline_md_N92, pipeline_md_N91, pipeline_md_N90,
         pipeline_md_N89, pipeline_md_N88, pipeline_md_N87, pipeline_md_N86,
         pipeline_md_N85, pipeline_md_N84, pipeline_md_N83, pipeline_md_N82,
         pipeline_md_N81, pipeline_md_N80, pipeline_md_N79, pipeline_md_N78,
         pipeline_md_N77, pipeline_md_N76, pipeline_md_N75, pipeline_md_N74,
         pipeline_md_N73, pipeline_md_N72, pipeline_md_N71, pipeline_md_N70,
         pipeline_md_N69, pipeline_md_N68, pipeline_md_N67, pipeline_md_N66,
         pipeline_md_N65, pipeline_md_N64, pipeline_md_N63, pipeline_md_N60,
         pipeline_md_N59, pipeline_md_N58, pipeline_md_N57, pipeline_md_N56,
         pipeline_md_N55, pipeline_md_N54, pipeline_md_N53, pipeline_md_N52,
         pipeline_md_N51, pipeline_md_N50, pipeline_md_N49, pipeline_md_N48,
         pipeline_md_N47, pipeline_md_N46, pipeline_md_N45, pipeline_md_N44,
         pipeline_md_N43, pipeline_md_N42, pipeline_md_N41, pipeline_md_N40,
         pipeline_md_N39, pipeline_md_N38, pipeline_md_N37, pipeline_md_N36,
         pipeline_md_N35, pipeline_md_N34, pipeline_md_N33, pipeline_md_N32,
         pipeline_md_N31, pipeline_md_N30, pipeline_md_N29, pipeline_md_N25,
         pipeline_md_N24, pipeline_md_N23, pipeline_md_N22, pipeline_md_N21,
         pipeline_csr_N2407, pipeline_csr_N2405, pipeline_csr_N2164,
         pipeline_csr_N2163, pipeline_csr_N2162, pipeline_csr_N2161,
         pipeline_csr_N2160, pipeline_csr_N2159, pipeline_csr_N2158,
         pipeline_csr_N2157, pipeline_csr_N2156, pipeline_csr_N2155,
         pipeline_csr_N2154, pipeline_csr_N2153, pipeline_csr_N2152,
         pipeline_csr_N2151, pipeline_csr_N2150, pipeline_csr_N2149,
         pipeline_csr_N2148, pipeline_csr_N2147, pipeline_csr_N2146,
         pipeline_csr_N2145, pipeline_csr_N2144, pipeline_csr_N2143,
         pipeline_csr_N2142, pipeline_csr_N2141, pipeline_csr_N2140,
         pipeline_csr_N2139, pipeline_csr_N2138, pipeline_csr_N2137,
         pipeline_csr_N2136, pipeline_csr_N2135, pipeline_csr_N2134,
         pipeline_csr_N2133, pipeline_csr_N2132, pipeline_csr_N2131,
         pipeline_csr_N2130, pipeline_csr_N2129, pipeline_csr_N2128,
         pipeline_csr_N2127, pipeline_csr_N2126, pipeline_csr_N2125,
         pipeline_csr_N2124, pipeline_csr_N2123, pipeline_csr_N2122,
         pipeline_csr_N2121, pipeline_csr_N2120, pipeline_csr_N2119,
         pipeline_csr_N2118, pipeline_csr_N2117, pipeline_csr_N2116,
         pipeline_csr_N2115, pipeline_csr_N2114, pipeline_csr_N2113,
         pipeline_csr_N2112, pipeline_csr_N2111, pipeline_csr_N2110,
         pipeline_csr_N2109, pipeline_csr_N2108, pipeline_csr_N2107,
         pipeline_csr_N2106, pipeline_csr_N2105, pipeline_csr_N2104,
         pipeline_csr_N2103, pipeline_csr_N2102, pipeline_csr_N2101,
         pipeline_csr_N2015, pipeline_csr_N2014, pipeline_csr_N2013,
         pipeline_csr_N2012, pipeline_csr_N2011, pipeline_csr_N2010,
         pipeline_csr_N2009, pipeline_csr_N2008, pipeline_csr_N2007,
         pipeline_csr_N2006, pipeline_csr_N2005, pipeline_csr_N2004,
         pipeline_csr_N2003, pipeline_csr_N2002, pipeline_csr_N2001,
         pipeline_csr_N2000, pipeline_csr_N1999, pipeline_csr_N1998,
         pipeline_csr_N1997, pipeline_csr_N1996, pipeline_csr_N1995,
         pipeline_csr_N1994, pipeline_csr_N1993, pipeline_csr_N1992,
         pipeline_csr_N1991, pipeline_csr_N1990, pipeline_csr_N1989,
         pipeline_csr_N1988, pipeline_csr_N1987, pipeline_csr_N1986,
         pipeline_csr_N1985, pipeline_csr_N1984, pipeline_csr_N1983,
         pipeline_csr_N1982, pipeline_csr_N1981, pipeline_csr_N1980,
         pipeline_csr_N1979, pipeline_csr_N1978, pipeline_csr_N1977,
         pipeline_csr_N1976, pipeline_csr_N1975, pipeline_csr_N1974,
         pipeline_csr_N1973, pipeline_csr_N1972, pipeline_csr_N1971,
         pipeline_csr_N1970, pipeline_csr_N1969, pipeline_csr_N1968,
         pipeline_csr_N1967, pipeline_csr_N1966, pipeline_csr_N1965,
         pipeline_csr_N1964, pipeline_csr_N1963, pipeline_csr_N1962,
         pipeline_csr_N1961, pipeline_csr_N1960, pipeline_csr_N1959,
         pipeline_csr_N1958, pipeline_csr_N1957, pipeline_csr_N1956,
         pipeline_csr_N1955, pipeline_csr_N1954, pipeline_csr_N1953,
         pipeline_csr_N1952, pipeline_csr_N1951, pipeline_csr_N1950,
         pipeline_csr_N1949, pipeline_csr_N1948, pipeline_csr_N1947,
         pipeline_csr_N1946, pipeline_csr_N1945, pipeline_csr_N1944,
         pipeline_csr_N1943, pipeline_csr_N1942, pipeline_csr_N1941,
         pipeline_csr_N1940, pipeline_csr_N1939, pipeline_csr_N1938,
         pipeline_csr_N1937, pipeline_csr_N1936, pipeline_csr_N1935,
         pipeline_csr_N1934, pipeline_csr_N1933, pipeline_csr_N1932,
         pipeline_csr_N1931, pipeline_csr_N1930, pipeline_csr_N1929,
         pipeline_csr_N1928, pipeline_csr_N1927, pipeline_csr_N1926,
         pipeline_csr_N1925, pipeline_csr_N1924, pipeline_csr_N1923,
         pipeline_csr_N1922, pipeline_csr_N1921, pipeline_csr_N1920,
         pipeline_csr_N1919, pipeline_csr_N1918, pipeline_csr_N1917,
         pipeline_csr_N1916, pipeline_csr_N1915, pipeline_csr_N1914,
         pipeline_csr_N1913, pipeline_csr_N1912, pipeline_csr_N1911,
         pipeline_csr_N1910, pipeline_csr_N1909, pipeline_csr_N1908,
         pipeline_csr_N1907, pipeline_csr_N1906, pipeline_csr_N1905,
         pipeline_csr_N1904, pipeline_csr_N1903, pipeline_csr_N1902,
         pipeline_csr_N1901, pipeline_csr_N1900, pipeline_csr_N1899,
         pipeline_csr_N1898, pipeline_csr_N1897, pipeline_csr_N1896,
         pipeline_csr_N1895, pipeline_csr_N1894, pipeline_csr_N1893,
         pipeline_csr_N1892, pipeline_csr_N1891, pipeline_csr_N1890,
         pipeline_csr_N1889, pipeline_csr_N1888, pipeline_csr_N903,
         pipeline_csr_N902, pipeline_csr_N901, pipeline_csr_N900,
         pipeline_csr_N899, pipeline_csr_N898, pipeline_csr_N897,
         pipeline_csr_N896, pipeline_csr_N895, pipeline_csr_N894,
         pipeline_csr_N893, pipeline_csr_N892, pipeline_csr_N891,
         pipeline_csr_N890, pipeline_csr_N889, pipeline_csr_N888,
         pipeline_csr_N887, pipeline_csr_N886, pipeline_csr_N885,
         pipeline_csr_N884, pipeline_csr_N883, pipeline_csr_N882,
         pipeline_csr_N881, pipeline_csr_N880, pipeline_csr_N879,
         pipeline_csr_N878, pipeline_csr_N877, pipeline_csr_N876,
         pipeline_csr_N875, pipeline_csr_N874, pipeline_csr_N873,
         pipeline_csr_N872, pipeline_csr_N871, pipeline_csr_N870,
         pipeline_csr_N869, pipeline_csr_N868, pipeline_csr_N867,
         pipeline_csr_N866, pipeline_csr_N865, pipeline_csr_N864,
         pipeline_csr_N863, pipeline_csr_N862, pipeline_csr_N861,
         pipeline_csr_N860, pipeline_csr_N859, pipeline_csr_N858,
         pipeline_csr_N857, pipeline_csr_N856, pipeline_csr_N855,
         pipeline_csr_N854, pipeline_csr_N853, pipeline_csr_N852,
         pipeline_csr_N851, pipeline_csr_N850, pipeline_csr_N849,
         pipeline_csr_N848, pipeline_csr_N847, pipeline_csr_N846,
         pipeline_csr_N845, pipeline_csr_N844, pipeline_csr_N843,
         pipeline_csr_N842, pipeline_csr_N841, pipeline_csr_N840,
         pipeline_csr_N839, pipeline_csr_N838, pipeline_csr_N837,
         pipeline_csr_N836, pipeline_csr_N835, pipeline_csr_N834,
         pipeline_csr_N833, pipeline_csr_N832, pipeline_csr_N831,
         pipeline_csr_N830, pipeline_csr_N829, pipeline_csr_N828,
         pipeline_csr_N827, pipeline_csr_N826, pipeline_csr_N825,
         pipeline_csr_N824, pipeline_csr_N823, pipeline_csr_N822,
         pipeline_csr_N821, pipeline_csr_N820, pipeline_csr_N819,
         pipeline_csr_N818, pipeline_csr_N817, pipeline_csr_N816,
         pipeline_csr_N815, pipeline_csr_N814, pipeline_csr_N813,
         pipeline_csr_N812, pipeline_csr_N811, pipeline_csr_N810,
         pipeline_csr_N809, pipeline_csr_N808, pipeline_csr_N807,
         pipeline_csr_N806, pipeline_csr_N805, pipeline_csr_N804,
         pipeline_csr_N803, pipeline_csr_N802, pipeline_csr_N801,
         pipeline_csr_N800, pipeline_csr_N799, pipeline_csr_N798,
         pipeline_csr_N797, pipeline_csr_N796, pipeline_csr_N795,
         pipeline_csr_N794, pipeline_csr_N793, pipeline_csr_N792,
         pipeline_csr_N791, pipeline_csr_N790, pipeline_csr_N789,
         pipeline_csr_N788, pipeline_csr_N787, pipeline_csr_N786,
         pipeline_csr_N785, pipeline_csr_N784, pipeline_csr_N783,
         pipeline_csr_N782, pipeline_csr_N781, pipeline_csr_N780,
         pipeline_csr_N779, pipeline_csr_N778, pipeline_csr_N777,
         pipeline_csr_N775, pipeline_csr_N774, pipeline_csr_N773,
         pipeline_csr_N772, pipeline_csr_N771, pipeline_csr_N770,
         pipeline_csr_N769, pipeline_csr_N768, pipeline_csr_N767,
         pipeline_csr_N766, pipeline_csr_N765, pipeline_csr_N764,
         pipeline_csr_N763, pipeline_csr_N762, pipeline_csr_N761,
         pipeline_csr_N760, pipeline_csr_N759, pipeline_csr_N758,
         pipeline_csr_N757, pipeline_csr_N756, pipeline_csr_N755,
         pipeline_csr_N754, pipeline_csr_N753, pipeline_csr_N752,
         pipeline_csr_N751, pipeline_csr_N750, pipeline_csr_N749,
         pipeline_csr_N748, pipeline_csr_N747, pipeline_csr_N746,
         pipeline_csr_N745, pipeline_csr_N744, pipeline_csr_N743,
         pipeline_csr_N742, pipeline_csr_N741, pipeline_csr_N740,
         pipeline_csr_N739, pipeline_csr_N738, pipeline_csr_N737,
         pipeline_csr_N736, pipeline_csr_N735, pipeline_csr_N734,
         pipeline_csr_N733, pipeline_csr_N732, pipeline_csr_N731,
         pipeline_csr_N730, pipeline_csr_N729, pipeline_csr_N728,
         pipeline_csr_N727, pipeline_csr_N726, pipeline_csr_N725,
         pipeline_csr_N724, pipeline_csr_N723, pipeline_csr_N722,
         pipeline_csr_N721, pipeline_csr_N720, pipeline_csr_N719,
         pipeline_csr_N718, pipeline_csr_N717, pipeline_csr_N716,
         pipeline_csr_N715, pipeline_csr_N714, pipeline_csr_N713,
         pipeline_csr_N712, pipeline_csr_N711, pipeline_csr_N710,
         pipeline_csr_N709, pipeline_csr_N708, pipeline_csr_N707,
         pipeline_csr_N706, pipeline_csr_N705, pipeline_csr_N704,
         pipeline_csr_N703, pipeline_csr_N702, pipeline_csr_N701,
         pipeline_csr_N700, pipeline_csr_N699, pipeline_csr_N698,
         pipeline_csr_N697, pipeline_csr_N696, pipeline_csr_N695,
         pipeline_csr_N694, pipeline_csr_N693, pipeline_csr_N692,
         pipeline_csr_N691, pipeline_csr_N690, pipeline_csr_N689,
         pipeline_csr_N688, pipeline_csr_N687, pipeline_csr_N686,
         pipeline_csr_N685, pipeline_csr_N684, pipeline_csr_N683,
         pipeline_csr_N682, pipeline_csr_N681, pipeline_csr_N680,
         pipeline_csr_N679, pipeline_csr_N678, pipeline_csr_N677,
         pipeline_csr_N676, pipeline_csr_N675, pipeline_csr_N674,
         pipeline_csr_N673, pipeline_csr_N672, pipeline_csr_N671,
         pipeline_csr_N670, pipeline_csr_N669, pipeline_csr_N668,
         pipeline_csr_N667, pipeline_csr_N666, pipeline_csr_N665,
         pipeline_csr_N664, pipeline_csr_N663, pipeline_csr_N662,
         pipeline_csr_N661, pipeline_csr_N660, pipeline_csr_N659,
         pipeline_csr_N658, pipeline_csr_N657, pipeline_csr_N656,
         pipeline_csr_N655, pipeline_csr_N654, pipeline_csr_N653,
         pipeline_csr_N652, pipeline_csr_N651, pipeline_csr_N650,
         pipeline_csr_N649, pipeline_csr_N648, pipeline_csr_to_host_3_,
         pipeline_csr_N332, pipeline_csr_N331, pipeline_csr_N330,
         pipeline_csr_N329, pipeline_csr_N328, pipeline_csr_N327,
         pipeline_csr_N326, pipeline_csr_N325, pipeline_csr_N324,
         pipeline_csr_N323, pipeline_csr_N322, pipeline_csr_N321,
         pipeline_csr_N320, pipeline_csr_N319, pipeline_csr_N318,
         pipeline_csr_N317, pipeline_csr_N316, pipeline_csr_N315,
         pipeline_csr_N314, pipeline_csr_N313, pipeline_csr_N312,
         pipeline_csr_N311, pipeline_csr_N310, pipeline_csr_N309,
         pipeline_csr_N308, pipeline_csr_N307, pipeline_csr_N306,
         pipeline_csr_N305, pipeline_csr_N304, pipeline_csr_N303,
         pipeline_csr_mip_3, pipeline_csr_mip_7_, pipeline_csr_N79,
         pipeline_csr_system_wen, pipeline_csr_priv_stack_0, n135, n136, n142,
         n143, n149, n150, n151, n152, n408, n410, n412, n414, n416, n418,
         n420, n422, n424, n426, n428, n430, n432, n434, n436, n438, n440,
         n442, n444, n446, n448, n450, n452, n454, n456, n458, n460, n462,
         n464, n466, n468, n470, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n594, n595, n596, n597, n598,
         n601, n602, n603, n636, n637, n638, n693, n700, n702, n713, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n780, n781,
         n784, n787, n789, n790, n791, n793, n799, n800, n898, n900, n902,
         n904, n906, n908, n910, n912, n914, n916, n918, n920, n922, n924,
         n926, n928, n930, n932, n934, n936, n938, n940, n942, n944, n946,
         n948, n950, n952, n954, n956, n958, n960, n962, n963, n964, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1087, n1088, n1091, n1092, n1095,
         n1096, n1099, n1100, n1103, n1104, n1107, n1108, n1111, n1112, n1115,
         n1116, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1153, n1154, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1195, n1196, n1197, n1198, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1226, n1228, n1229, n1231, n1238, n1243, n1251, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1319, n1384, n1385,
         n1387, n1389, n1418, n1420, n1422, n1423, n1430, n1435, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1447, n1448, n1478, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1549, n1558, n1562,
         n1905, n1907, n1909, n1911, n1915, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n3683, n3689, n3704, n3711, n3715, n3718, n3721, n3724, n3727, n3730,
         n3733, n3736, n3739, n3742, n3745, n3748, n3751, n3754, n3757, n3760,
         n3785, n4130, n4147, n4148, n4149, n4150, n4151, n4184, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4229, n4230, n4231, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9342, n9344, n9346, n9348,
         n9350, n9352, n9354, n9356, n9358, n9360, n9362, n9364, n9366, n9368,
         n9370, n9372, n9374, n9376, n9378, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5;
  wire   [2:0] pipeline_dmem_type_WB;
  wire   [31:0] pipeline_alu_out_WB;
  wire   [31:0] pipeline_md_resp_result;
  wire   [30:0] pipeline_alu_src_b;
  wire   [31:0] pipeline_rs2_data_bypassed;
  wire   [30:0] pipeline_alu_src_a;
  wire   [31:2] pipeline_handler_PC;
  wire   [31:0] pipeline_PC_DX;
  wire   [31:0] pipeline_rs1_data_bypassed;
  wire   [2:1] pipeline_reg_to_wr_WB;
  wire   [30:0] pipeline_inst_DX;
  wire   [3:0] pipeline_ctrl_prev_ex_code_WB;
  wire   [19:1] pipeline_PCmux_offset;
  wire   [31:0] pipeline_PCmux_base;
  wire   [1023:0] pipeline_regfile_data;
  wire   [63:0] pipeline_md_result_muxed;
  wire   [1:0] pipeline_md_out_sel;
  wire   [63:0] pipeline_md_b;
  wire   [62:0] pipeline_md_a;
  wire   [62:32] pipeline_md_result;
  wire   [1:0] pipeline_md_state;
  wire   [31:6] pipeline_csr_mscratch;
  wire   [63:0] pipeline_csr_instret_full;
  wire   [63:0] pipeline_csr_time_full;
  wire   [63:0] pipeline_csr_cycle_full;
  wire   [31:0] pipeline_csr_from_host;
  wire   [3:0] pipeline_csr_mbadaddr;
  wire   [63:0] pipeline_csr_mtime_full;
  wire   [31:0] pipeline_csr_mtimecmp;
  wire   [31:7] pipeline_csr_mie;
  wire   [6:0] pipeline_csr_mtvec;
  assign dmem_hsize[2] = 1'b0;
  assign dmem_htrans[0] = 1'b0;
  assign htif_pcr_resp_data[63] = 1'b0;
  assign htif_pcr_resp_data[62] = 1'b0;
  assign htif_pcr_resp_data[61] = 1'b0;
  assign htif_pcr_resp_data[60] = 1'b0;
  assign htif_pcr_resp_data[59] = 1'b0;
  assign htif_pcr_resp_data[58] = 1'b0;
  assign htif_pcr_resp_data[57] = 1'b0;
  assign htif_pcr_resp_data[56] = 1'b0;
  assign htif_pcr_resp_data[55] = 1'b0;
  assign htif_pcr_resp_data[54] = 1'b0;
  assign htif_pcr_resp_data[53] = 1'b0;
  assign htif_pcr_resp_data[52] = 1'b0;
  assign htif_pcr_resp_data[51] = 1'b0;
  assign htif_pcr_resp_data[50] = 1'b0;
  assign htif_pcr_resp_data[49] = 1'b0;
  assign htif_pcr_resp_data[48] = 1'b0;
  assign htif_pcr_resp_data[47] = 1'b0;
  assign htif_pcr_resp_data[46] = 1'b0;
  assign htif_pcr_resp_data[45] = 1'b0;
  assign htif_pcr_resp_data[44] = 1'b0;
  assign htif_pcr_resp_data[43] = 1'b0;
  assign htif_pcr_resp_data[42] = 1'b0;
  assign htif_pcr_resp_data[41] = 1'b0;
  assign htif_pcr_resp_data[40] = 1'b0;
  assign htif_pcr_resp_data[39] = 1'b0;
  assign htif_pcr_resp_data[38] = 1'b0;
  assign htif_pcr_resp_data[37] = 1'b0;
  assign htif_pcr_resp_data[36] = 1'b0;
  assign htif_pcr_resp_data[35] = 1'b0;
  assign htif_pcr_resp_data[34] = 1'b0;
  assign htif_pcr_resp_data[33] = 1'b0;
  assign htif_pcr_resp_data[32] = 1'b0;
  assign htif_debug_stats_pcr = 1'b0;
  assign htif_ipi_req_data = 1'b0;
  assign htif_ipi_req_valid = 1'b0;
  assign dmem_hprot[3] = 1'b0;
  assign dmem_hprot[2] = 1'b0;
  assign dmem_hprot[1] = 1'b0;
  assign dmem_hprot[0] = 1'b0;
  assign dmem_hmastlock = 1'b0;
  assign dmem_hburst[2] = 1'b0;
  assign dmem_hburst[1] = 1'b0;
  assign dmem_hburst[0] = 1'b0;
  assign imem_hwdata[31] = 1'b0;
  assign imem_hwdata[30] = 1'b0;
  assign imem_hwdata[29] = 1'b0;
  assign imem_hwdata[28] = 1'b0;
  assign imem_hwdata[27] = 1'b0;
  assign imem_hwdata[26] = 1'b0;
  assign imem_hwdata[25] = 1'b0;
  assign imem_hwdata[24] = 1'b0;
  assign imem_hwdata[23] = 1'b0;
  assign imem_hwdata[22] = 1'b0;
  assign imem_hwdata[21] = 1'b0;
  assign imem_hwdata[20] = 1'b0;
  assign imem_hwdata[19] = 1'b0;
  assign imem_hwdata[18] = 1'b0;
  assign imem_hwdata[17] = 1'b0;
  assign imem_hwdata[16] = 1'b0;
  assign imem_hwdata[15] = 1'b0;
  assign imem_hwdata[14] = 1'b0;
  assign imem_hwdata[13] = 1'b0;
  assign imem_hwdata[12] = 1'b0;
  assign imem_hwdata[11] = 1'b0;
  assign imem_hwdata[10] = 1'b0;
  assign imem_hwdata[9] = 1'b0;
  assign imem_hwdata[8] = 1'b0;
  assign imem_hwdata[7] = 1'b0;
  assign imem_hwdata[6] = 1'b0;
  assign imem_hwdata[5] = 1'b0;
  assign imem_hwdata[4] = 1'b0;
  assign imem_hwdata[3] = 1'b0;
  assign imem_hwdata[2] = 1'b0;
  assign imem_hwdata[1] = 1'b0;
  assign imem_hwdata[0] = 1'b0;
  assign imem_htrans[1] = 1'b1;
  assign imem_htrans[0] = 1'b0;
  assign imem_hprot[3] = 1'b0;
  assign imem_hprot[2] = 1'b0;
  assign imem_hprot[1] = 1'b0;
  assign imem_hprot[0] = 1'b0;
  assign imem_hmastlock = 1'b0;
  assign imem_hburst[2] = 1'b0;
  assign imem_hburst[1] = 1'b0;
  assign imem_hburst[0] = 1'b0;
  assign imem_hsize[2] = 1'b0;
  assign imem_hsize[1] = 1'b1;
  assign imem_hsize[0] = 1'b0;
  assign imem_hwrite = 1'b0;
  assign htif_ipi_resp_ready = 1'b1;

  vscale_core_DW_cmp_0 pipeline_md_gte_63 

  INV_X4 vscale_core_DW_cmp_0_U313 ( .A(vscale_core_DW_cmp_0n545), .ZN(vscale_core_DW_cmp_0n446) );
  INV_X4 vscale_core_DW_cmp_0_U314 ( .A(vscale_core_DW_cmp_0n580), .ZN(vscale_core_DW_cmp_0n447) );
  INV_X4 vscale_core_DW_cmp_0_U315 ( .A(pipeline_md_b[31]), .ZN(vscale_core_DW_cmp_0n448) );
  INV_X4 vscale_core_DW_cmp_0_U316 ( .A(pipeline_md_b[29]), .ZN(vscale_core_DW_cmp_0n449) );
  INV_X4 vscale_core_DW_cmp_0_U317 ( .A(vscale_core_DW_cmp_0n573), .ZN(vscale_core_DW_cmp_0n450) );
  INV_X4 vscale_core_DW_cmp_0_U318 ( .A(pipeline_md_b[27]), .ZN(vscale_core_DW_cmp_0n451) );
  INV_X4 vscale_core_DW_cmp_0_U319 ( .A(pipeline_md_b[25]), .ZN(vscale_core_DW_cmp_0n452) );
  INV_X4 vscale_core_DW_cmp_0_U320 ( .A(vscale_core_DW_cmp_0n578), .ZN(vscale_core_DW_cmp_0n453) );
  INV_X4 vscale_core_DW_cmp_0_U321 ( .A(pipeline_md_b[23]), .ZN(vscale_core_DW_cmp_0n454) );
  INV_X4 vscale_core_DW_cmp_0_U322 ( .A(pipeline_md_b[21]), .ZN(vscale_core_DW_cmp_0n455) );
  INV_X4 vscale_core_DW_cmp_0_U323 ( .A(vscale_core_DW_cmp_0n557), .ZN(vscale_core_DW_cmp_0n456) );
  INV_X4 vscale_core_DW_cmp_0_U324 ( .A(pipeline_md_b[19]), .ZN(vscale_core_DW_cmp_0n457) );
  INV_X4 vscale_core_DW_cmp_0_U325 ( .A(pipeline_md_b[17]), .ZN(vscale_core_DW_cmp_0n458) );
  INV_X4 vscale_core_DW_cmp_0_U326 ( .A(vscale_core_DW_cmp_0n604), .ZN(vscale_core_DW_cmp_0n459) );
  INV_X4 vscale_core_DW_cmp_0_U327 ( .A(vscale_core_DW_cmp_0n618), .ZN(vscale_core_DW_cmp_0n460) );
  INV_X4 vscale_core_DW_cmp_0_U328 ( .A(pipeline_md_b[15]), .ZN(vscale_core_DW_cmp_0n461) );
  INV_X4 vscale_core_DW_cmp_0_U329 ( .A(pipeline_md_b[13]), .ZN(vscale_core_DW_cmp_0n462) );
  INV_X4 vscale_core_DW_cmp_0_U330 ( .A(vscale_core_DW_cmp_0n603), .ZN(vscale_core_DW_cmp_0n463) );
  INV_X4 vscale_core_DW_cmp_0_U331 ( .A(pipeline_md_b[11]), .ZN(vscale_core_DW_cmp_0n464) );
  INV_X4 vscale_core_DW_cmp_0_U332 ( .A(pipeline_md_b[9]), .ZN(vscale_core_DW_cmp_0n465) );
  INV_X4 vscale_core_DW_cmp_0_U333 ( .A(vscale_core_DW_cmp_0n591), .ZN(vscale_core_DW_cmp_0n466) );
  INV_X4 vscale_core_DW_cmp_0_U334 ( .A(pipeline_md_b[7]), .ZN(vscale_core_DW_cmp_0n467) );
  INV_X4 vscale_core_DW_cmp_0_U335 ( .A(pipeline_md_b[4]), .ZN(vscale_core_DW_cmp_0n468) );
  INV_X4 vscale_core_DW_cmp_0_U336 ( .A(vscale_core_DW_cmp_0n597), .ZN(vscale_core_DW_cmp_0n469) );
  INV_X4 vscale_core_DW_cmp_0_U337 ( .A(pipeline_md_b[3]), .ZN(vscale_core_DW_cmp_0n470) );
  INV_X4 vscale_core_DW_cmp_0_U338 ( .A(pipeline_md_b[1]), .ZN(vscale_core_DW_cmp_0n471) );
  INV_X4 vscale_core_DW_cmp_0_U339 ( .A(vscale_core_DW_cmp_0n539), .ZN(vscale_core_DW_cmp_0n472) );
  INV_X4 vscale_core_DW_cmp_0_U340 ( .A(vscale_core_DW_cmp_0n623), .ZN(vscale_core_DW_cmp_0n473) );
  INV_X4 vscale_core_DW_cmp_0_U341 ( .A(vscale_core_DW_cmp_0n689), .ZN(vscale_core_DW_cmp_0n474) );
  INV_X4 vscale_core_DW_cmp_0_U342 ( .A(n10233), .ZN(vscale_core_DW_cmp_0n475) );
  INV_X4 vscale_core_DW_cmp_0_U343 ( .A(pipeline_md_a[30]), .ZN(vscale_core_DW_cmp_0n476) );
  INV_X4 vscale_core_DW_cmp_0_U344 ( .A(pipeline_md_a[32]), .ZN(vscale_core_DW_cmp_0n477) );
  INV_X4 vscale_core_DW_cmp_0_U345 ( .A(vscale_core_DW_cmp_0n535), .ZN(vscale_core_DW_cmp_0n478) );
  INV_X4 vscale_core_DW_cmp_0_U346 ( .A(pipeline_md_a[34]), .ZN(vscale_core_DW_cmp_0n479) );
  INV_X4 vscale_core_DW_cmp_0_U347 ( .A(pipeline_md_a[36]), .ZN(vscale_core_DW_cmp_0n480) );
  INV_X4 vscale_core_DW_cmp_0_U348 ( .A(vscale_core_DW_cmp_0n671), .ZN(vscale_core_DW_cmp_0n481) );
  INV_X4 vscale_core_DW_cmp_0_U349 ( .A(pipeline_md_a[38]), .ZN(vscale_core_DW_cmp_0n482) );
  INV_X4 vscale_core_DW_cmp_0_U350 ( .A(vscale_core_DW_cmp_0n537), .ZN(vscale_core_DW_cmp_0n483) );
  INV_X4 vscale_core_DW_cmp_0_U351 ( .A(pipeline_md_a[40]), .ZN(vscale_core_DW_cmp_0n484) );
  INV_X4 vscale_core_DW_cmp_0_U352 ( .A(vscale_core_DW_cmp_0n657), .ZN(vscale_core_DW_cmp_0n485) );
  INV_X4 vscale_core_DW_cmp_0_U353 ( .A(pipeline_md_a[42]), .ZN(vscale_core_DW_cmp_0n486) );
  INV_X4 vscale_core_DW_cmp_0_U354 ( .A(pipeline_md_a[44]), .ZN(vscale_core_DW_cmp_0n487) );
  INV_X4 vscale_core_DW_cmp_0_U355 ( .A(vscale_core_DW_cmp_0n685), .ZN(vscale_core_DW_cmp_0n488) );
  INV_X4 vscale_core_DW_cmp_0_U356 ( .A(pipeline_md_a[46]), .ZN(vscale_core_DW_cmp_0n489) );
  INV_X4 vscale_core_DW_cmp_0_U357 ( .A(pipeline_md_a[48]), .ZN(vscale_core_DW_cmp_0n490) );
  INV_X4 vscale_core_DW_cmp_0_U358 ( .A(vscale_core_DW_cmp_0n635), .ZN(vscale_core_DW_cmp_0n491) );
  INV_X4 vscale_core_DW_cmp_0_U359 ( .A(pipeline_md_a[50]), .ZN(vscale_core_DW_cmp_0n492) );
  INV_X4 vscale_core_DW_cmp_0_U360 ( .A(pipeline_md_a[52]), .ZN(vscale_core_DW_cmp_0n493) );
  INV_X4 vscale_core_DW_cmp_0_U361 ( .A(vscale_core_DW_cmp_0n687), .ZN(vscale_core_DW_cmp_0n494) );
  INV_X4 vscale_core_DW_cmp_0_U362 ( .A(pipeline_md_a[54]), .ZN(vscale_core_DW_cmp_0n495) );
  INV_X4 vscale_core_DW_cmp_0_U363 ( .A(pipeline_md_a[56]), .ZN(vscale_core_DW_cmp_0n496) );
  INV_X4 vscale_core_DW_cmp_0_U364 ( .A(vscale_core_DW_cmp_0n645), .ZN(vscale_core_DW_cmp_0n497) );
  INV_X4 vscale_core_DW_cmp_0_U365 ( .A(pipeline_md_a[58]), .ZN(vscale_core_DW_cmp_0n498) );
  INV_X4 vscale_core_DW_cmp_0_U366 ( .A(pipeline_md_a[61]), .ZN(vscale_core_DW_cmp_0n499) );
  INV_X4 vscale_core_DW_cmp_0_U367 ( .A(pipeline_md_a[5]), .ZN(vscale_core_DW_cmp_0n500) );
  INV_X4 vscale_core_DW_cmp_0_U368 ( .A(pipeline_md_a[1]), .ZN(vscale_core_DW_cmp_0n501) );
  INV_X4 vscale_core_DW_cmp_0_U369 ( .A(pipeline_md_a[2]), .ZN(vscale_core_DW_cmp_0n502) );
  INV_X4 vscale_core_DW_cmp_0_U370 ( .A(pipeline_md_a[6]), .ZN(vscale_core_DW_cmp_0n503) );
  INV_X4 vscale_core_DW_cmp_0_U371 ( .A(pipeline_md_a[8]), .ZN(vscale_core_DW_cmp_0n504) );
  INV_X4 vscale_core_DW_cmp_0_U372 ( .A(pipeline_md_a[10]), .ZN(vscale_core_DW_cmp_0n505) );
  INV_X4 vscale_core_DW_cmp_0_U373 ( .A(pipeline_md_a[12]), .ZN(vscale_core_DW_cmp_0n506) );
  INV_X4 vscale_core_DW_cmp_0_U374 ( .A(pipeline_md_a[14]), .ZN(vscale_core_DW_cmp_0n507) );
  INV_X4 vscale_core_DW_cmp_0_U375 ( .A(pipeline_md_a[16]), .ZN(vscale_core_DW_cmp_0n508) );
  INV_X4 vscale_core_DW_cmp_0_U376 ( .A(pipeline_md_a[18]), .ZN(vscale_core_DW_cmp_0n509) );
  INV_X4 vscale_core_DW_cmp_0_U377 ( .A(pipeline_md_a[20]), .ZN(vscale_core_DW_cmp_0n510) );
  INV_X4 vscale_core_DW_cmp_0_U378 ( .A(pipeline_md_b[60]), .ZN(vscale_core_DW_cmp_0n511) );
  INV_X4 vscale_core_DW_cmp_0_U379 ( .A(pipeline_md_b[59]), .ZN(vscale_core_DW_cmp_0n512) );
  INV_X4 vscale_core_DW_cmp_0_U380 ( .A(pipeline_md_b[57]), .ZN(vscale_core_DW_cmp_0n513) );
  INV_X4 vscale_core_DW_cmp_0_U381 ( .A(pipeline_md_b[55]), .ZN(vscale_core_DW_cmp_0n514) );
  INV_X4 vscale_core_DW_cmp_0_U382 ( .A(pipeline_md_b[53]), .ZN(vscale_core_DW_cmp_0n515) );
  INV_X4 vscale_core_DW_cmp_0_U383 ( .A(pipeline_md_b[51]), .ZN(vscale_core_DW_cmp_0n516) );
  INV_X4 vscale_core_DW_cmp_0_U384 ( .A(pipeline_md_b[49]), .ZN(vscale_core_DW_cmp_0n517) );
  INV_X4 vscale_core_DW_cmp_0_U385 ( .A(pipeline_md_b[47]), .ZN(vscale_core_DW_cmp_0n518) );
  INV_X4 vscale_core_DW_cmp_0_U386 ( .A(pipeline_md_b[45]), .ZN(vscale_core_DW_cmp_0n519) );
  INV_X4 vscale_core_DW_cmp_0_U387 ( .A(pipeline_md_b[43]), .ZN(vscale_core_DW_cmp_0n520) );
  INV_X4 vscale_core_DW_cmp_0_U388 ( .A(pipeline_md_b[41]), .ZN(vscale_core_DW_cmp_0n521) );
  INV_X4 vscale_core_DW_cmp_0_U389 ( .A(pipeline_md_b[39]), .ZN(vscale_core_DW_cmp_0n522) );
  INV_X4 vscale_core_DW_cmp_0_U390 ( .A(pipeline_md_b[37]), .ZN(vscale_core_DW_cmp_0n523) );
  INV_X4 vscale_core_DW_cmp_0_U391 ( .A(pipeline_md_b[35]), .ZN(vscale_core_DW_cmp_0n524) );
  INV_X4 vscale_core_DW_cmp_0_U392 ( .A(pipeline_md_b[33]), .ZN(vscale_core_DW_cmp_0n525) );
  INV_X4 vscale_core_DW_cmp_0_U393 ( .A(pipeline_md_a[22]), .ZN(vscale_core_DW_cmp_0n526) );
  INV_X4 vscale_core_DW_cmp_0_U394 ( .A(pipeline_md_a[24]), .ZN(vscale_core_DW_cmp_0n527) );
  INV_X4 vscale_core_DW_cmp_0_U395 ( .A(pipeline_md_a[26]), .ZN(vscale_core_DW_cmp_0n528) );
  INV_X4 vscale_core_DW_cmp_0_U396 ( .A(pipeline_md_a[28]), .ZN(vscale_core_DW_cmp_0n529) );
  INV_X4 vscale_core_DW_cmp_0_U397 ( .A(pipeline_md_a[62]), .ZN(vscale_core_DW_cmp_0n530) );
  OAI22_X1 vscale_core_DW_cmp_0_U398 ( .A1(vscale_core_DW_cmp_0n531), .A2(vscale_core_DW_cmp_0n532), .B1(vscale_core_DW_cmp_0n533), .B2(vscale_core_DW_cmp_0n531), .ZN(pipeline_md_a_geq)
         );
  NOR4_X1 vscale_core_DW_cmp_0_U399 ( .A1(vscale_core_DW_cmp_0n534), .A2(vscale_core_DW_cmp_0n535), .A3(vscale_core_DW_cmp_0n536), .A4(vscale_core_DW_cmp_0n537), .ZN(vscale_core_DW_cmp_0n533) );
  OAI211_X1 vscale_core_DW_cmp_0_U400 ( .C1(pipeline_md_b[32]), .C2(vscale_core_DW_cmp_0n477), .A(vscale_core_DW_cmp_0n538), .B(vscale_core_DW_cmp_0n539), .ZN(vscale_core_DW_cmp_0n534) );
  OAI21_X1 vscale_core_DW_cmp_0_U401 ( .B1(vscale_core_DW_cmp_0n540), .B2(vscale_core_DW_cmp_0n541), .A(vscale_core_DW_cmp_0n542), .ZN(vscale_core_DW_cmp_0n532) );
  OAI22_X1 vscale_core_DW_cmp_0_U402 ( .A1(vscale_core_DW_cmp_0n543), .A2(vscale_core_DW_cmp_0n544), .B1(vscale_core_DW_cmp_0n446), .B2(vscale_core_DW_cmp_0n543), .ZN(vscale_core_DW_cmp_0n542) );
  OAI21_X1 vscale_core_DW_cmp_0_U403 ( .B1(vscale_core_DW_cmp_0n546), .B2(vscale_core_DW_cmp_0n547), .A(vscale_core_DW_cmp_0n548), .ZN(vscale_core_DW_cmp_0n544) );
  OAI22_X1 vscale_core_DW_cmp_0_U404 ( .A1(vscale_core_DW_cmp_0n549), .A2(vscale_core_DW_cmp_0n550), .B1(vscale_core_DW_cmp_0n453), .B2(vscale_core_DW_cmp_0n549), .ZN(vscale_core_DW_cmp_0n548) );
  OAI21_X1 vscale_core_DW_cmp_0_U405 ( .B1(pipeline_md_a[21]), .B2(vscale_core_DW_cmp_0n455), .A(vscale_core_DW_cmp_0n551), .ZN(vscale_core_DW_cmp_0n550) );
  NAND3_X1 vscale_core_DW_cmp_0_U406 ( .A1(vscale_core_DW_cmp_0n552), .A2(vscale_core_DW_cmp_0n510), .A3(pipeline_md_b[20]), .ZN(vscale_core_DW_cmp_0n551) );
  OAI21_X1 vscale_core_DW_cmp_0_U407 ( .B1(pipeline_md_a[23]), .B2(vscale_core_DW_cmp_0n454), .A(vscale_core_DW_cmp_0n553), .ZN(vscale_core_DW_cmp_0n549) );
  NAND3_X1 vscale_core_DW_cmp_0_U408 ( .A1(vscale_core_DW_cmp_0n554), .A2(vscale_core_DW_cmp_0n526), .A3(pipeline_md_b[22]), .ZN(vscale_core_DW_cmp_0n553) );
  OAI22_X1 vscale_core_DW_cmp_0_U409 ( .A1(vscale_core_DW_cmp_0n555), .A2(vscale_core_DW_cmp_0n556), .B1(vscale_core_DW_cmp_0n456), .B2(vscale_core_DW_cmp_0n555), .ZN(vscale_core_DW_cmp_0n547) );
  OAI21_X1 vscale_core_DW_cmp_0_U410 ( .B1(pipeline_md_a[17]), .B2(vscale_core_DW_cmp_0n458), .A(vscale_core_DW_cmp_0n558), .ZN(vscale_core_DW_cmp_0n556) );
  NAND3_X1 vscale_core_DW_cmp_0_U411 ( .A1(vscale_core_DW_cmp_0n559), .A2(vscale_core_DW_cmp_0n508), .A3(pipeline_md_b[16]), .ZN(vscale_core_DW_cmp_0n558) );
  OAI21_X1 vscale_core_DW_cmp_0_U412 ( .B1(pipeline_md_a[19]), .B2(vscale_core_DW_cmp_0n457), .A(vscale_core_DW_cmp_0n560), .ZN(vscale_core_DW_cmp_0n555) );
  NAND3_X1 vscale_core_DW_cmp_0_U413 ( .A1(vscale_core_DW_cmp_0n561), .A2(vscale_core_DW_cmp_0n509), .A3(pipeline_md_b[18]), .ZN(vscale_core_DW_cmp_0n560) );
  OAI21_X1 vscale_core_DW_cmp_0_U414 ( .B1(vscale_core_DW_cmp_0n562), .B2(vscale_core_DW_cmp_0n563), .A(vscale_core_DW_cmp_0n564), .ZN(vscale_core_DW_cmp_0n543) );
  OAI22_X1 vscale_core_DW_cmp_0_U415 ( .A1(vscale_core_DW_cmp_0n565), .A2(vscale_core_DW_cmp_0n566), .B1(vscale_core_DW_cmp_0n447), .B2(vscale_core_DW_cmp_0n565), .ZN(vscale_core_DW_cmp_0n564) );
  OAI21_X1 vscale_core_DW_cmp_0_U416 ( .B1(pipeline_md_a[29]), .B2(vscale_core_DW_cmp_0n449), .A(vscale_core_DW_cmp_0n567), .ZN(vscale_core_DW_cmp_0n566) );
  NAND3_X1 vscale_core_DW_cmp_0_U417 ( .A1(vscale_core_DW_cmp_0n568), .A2(vscale_core_DW_cmp_0n529), .A3(pipeline_md_b[28]), .ZN(vscale_core_DW_cmp_0n567) );
  OAI21_X1 vscale_core_DW_cmp_0_U418 ( .B1(pipeline_md_a[31]), .B2(vscale_core_DW_cmp_0n448), .A(vscale_core_DW_cmp_0n569), .ZN(vscale_core_DW_cmp_0n565) );
  NAND3_X1 vscale_core_DW_cmp_0_U419 ( .A1(vscale_core_DW_cmp_0n570), .A2(vscale_core_DW_cmp_0n476), .A3(pipeline_md_b[30]), .ZN(vscale_core_DW_cmp_0n569) );
  OAI22_X1 vscale_core_DW_cmp_0_U420 ( .A1(vscale_core_DW_cmp_0n571), .A2(vscale_core_DW_cmp_0n572), .B1(vscale_core_DW_cmp_0n450), .B2(vscale_core_DW_cmp_0n571), .ZN(vscale_core_DW_cmp_0n563) );
  OAI21_X1 vscale_core_DW_cmp_0_U421 ( .B1(pipeline_md_a[25]), .B2(vscale_core_DW_cmp_0n452), .A(vscale_core_DW_cmp_0n574), .ZN(vscale_core_DW_cmp_0n572) );
  NAND3_X1 vscale_core_DW_cmp_0_U422 ( .A1(vscale_core_DW_cmp_0n575), .A2(vscale_core_DW_cmp_0n527), .A3(pipeline_md_b[24]), .ZN(vscale_core_DW_cmp_0n574) );
  OAI21_X1 vscale_core_DW_cmp_0_U423 ( .B1(pipeline_md_a[27]), .B2(vscale_core_DW_cmp_0n451), .A(vscale_core_DW_cmp_0n576), .ZN(vscale_core_DW_cmp_0n571) );
  NAND3_X1 vscale_core_DW_cmp_0_U424 ( .A1(vscale_core_DW_cmp_0n577), .A2(vscale_core_DW_cmp_0n528), .A3(pipeline_md_b[26]), .ZN(vscale_core_DW_cmp_0n576) );
  OR3_X1 vscale_core_DW_cmp_0_U425 ( .A1(vscale_core_DW_cmp_0n545), .A2(vscale_core_DW_cmp_0n546), .A3(vscale_core_DW_cmp_0n557), .ZN(vscale_core_DW_cmp_0n541) );
  OAI21_X1 vscale_core_DW_cmp_0_U426 ( .B1(pipeline_md_b[18]), .B2(vscale_core_DW_cmp_0n509), .A(vscale_core_DW_cmp_0n561), .ZN(vscale_core_DW_cmp_0n557) );
  NAND2_X1 vscale_core_DW_cmp_0_U427 ( .A1(pipeline_md_a[19]), .A2(vscale_core_DW_cmp_0n457), .ZN(vscale_core_DW_cmp_0n561) );
  OAI211_X1 vscale_core_DW_cmp_0_U428 ( .C1(pipeline_md_b[20]), .C2(vscale_core_DW_cmp_0n510), .A(vscale_core_DW_cmp_0n552), .B(vscale_core_DW_cmp_0n453), .ZN(vscale_core_DW_cmp_0n546) );
  OAI21_X1 vscale_core_DW_cmp_0_U429 ( .B1(pipeline_md_b[22]), .B2(vscale_core_DW_cmp_0n526), .A(vscale_core_DW_cmp_0n554), .ZN(vscale_core_DW_cmp_0n578) );
  NAND2_X1 vscale_core_DW_cmp_0_U430 ( .A1(pipeline_md_a[23]), .A2(vscale_core_DW_cmp_0n454), .ZN(vscale_core_DW_cmp_0n554) );
  NAND2_X1 vscale_core_DW_cmp_0_U431 ( .A1(pipeline_md_a[21]), .A2(vscale_core_DW_cmp_0n455), .ZN(vscale_core_DW_cmp_0n552) );
  OAI211_X1 vscale_core_DW_cmp_0_U432 ( .C1(pipeline_md_b[24]), .C2(vscale_core_DW_cmp_0n527), .A(vscale_core_DW_cmp_0n575), .B(vscale_core_DW_cmp_0n579), .ZN(vscale_core_DW_cmp_0n545) );
  NOR2_X1 vscale_core_DW_cmp_0_U433 ( .A1(vscale_core_DW_cmp_0n562), .A2(vscale_core_DW_cmp_0n573), .ZN(vscale_core_DW_cmp_0n579) );
  OAI21_X1 vscale_core_DW_cmp_0_U434 ( .B1(pipeline_md_b[26]), .B2(vscale_core_DW_cmp_0n528), .A(vscale_core_DW_cmp_0n577), .ZN(vscale_core_DW_cmp_0n573) );
  NAND2_X1 vscale_core_DW_cmp_0_U435 ( .A1(pipeline_md_a[27]), .A2(vscale_core_DW_cmp_0n451), .ZN(vscale_core_DW_cmp_0n577) );
  OAI211_X1 vscale_core_DW_cmp_0_U436 ( .C1(pipeline_md_b[28]), .C2(vscale_core_DW_cmp_0n529), .A(vscale_core_DW_cmp_0n568), .B(vscale_core_DW_cmp_0n447), .ZN(vscale_core_DW_cmp_0n562) );
  OAI21_X1 vscale_core_DW_cmp_0_U437 ( .B1(pipeline_md_b[30]), .B2(vscale_core_DW_cmp_0n476), .A(vscale_core_DW_cmp_0n570), .ZN(vscale_core_DW_cmp_0n580) );
  NAND2_X1 vscale_core_DW_cmp_0_U438 ( .A1(pipeline_md_a[31]), .A2(vscale_core_DW_cmp_0n448), .ZN(vscale_core_DW_cmp_0n570) );
  NAND2_X1 vscale_core_DW_cmp_0_U439 ( .A1(pipeline_md_a[29]), .A2(vscale_core_DW_cmp_0n449), .ZN(vscale_core_DW_cmp_0n568) );
  NAND2_X1 vscale_core_DW_cmp_0_U440 ( .A1(pipeline_md_a[25]), .A2(vscale_core_DW_cmp_0n452), .ZN(vscale_core_DW_cmp_0n575) );
  OAI211_X1 vscale_core_DW_cmp_0_U441 ( .C1(pipeline_md_b[16]), .C2(vscale_core_DW_cmp_0n508), .A(vscale_core_DW_cmp_0n559), .B(vscale_core_DW_cmp_0n581), .ZN(vscale_core_DW_cmp_0n540) );
  AOI22_X1 vscale_core_DW_cmp_0_U442 ( .A1(vscale_core_DW_cmp_0n459), .A2(vscale_core_DW_cmp_0n582), .B1(vscale_core_DW_cmp_0n583), .B2(vscale_core_DW_cmp_0n459), .ZN(vscale_core_DW_cmp_0n581) );
  AOI21_X1 vscale_core_DW_cmp_0_U443 ( .B1(vscale_core_DW_cmp_0n584), .B2(vscale_core_DW_cmp_0n585), .A(vscale_core_DW_cmp_0n586), .ZN(vscale_core_DW_cmp_0n583) );
  AOI22_X1 vscale_core_DW_cmp_0_U444 ( .A1(vscale_core_DW_cmp_0n466), .A2(vscale_core_DW_cmp_0n587), .B1(vscale_core_DW_cmp_0n588), .B2(vscale_core_DW_cmp_0n466), .ZN(vscale_core_DW_cmp_0n586) );
  AOI22_X1 vscale_core_DW_cmp_0_U445 ( .A1(pipeline_md_b[5]), .A2(vscale_core_DW_cmp_0n500), .B1(vscale_core_DW_cmp_0n589), .B2(pipeline_md_b[4]), .ZN(vscale_core_DW_cmp_0n588) );
  NOR2_X1 vscale_core_DW_cmp_0_U446 ( .A1(pipeline_md_a[4]), .A2(vscale_core_DW_cmp_0n590), .ZN(vscale_core_DW_cmp_0n589) );
  OAI21_X1 vscale_core_DW_cmp_0_U447 ( .B1(pipeline_md_a[7]), .B2(vscale_core_DW_cmp_0n467), .A(vscale_core_DW_cmp_0n592), .ZN(vscale_core_DW_cmp_0n591) );
  NAND3_X1 vscale_core_DW_cmp_0_U448 ( .A1(vscale_core_DW_cmp_0n593), .A2(vscale_core_DW_cmp_0n503), .A3(pipeline_md_b[6]), .ZN(vscale_core_DW_cmp_0n592) );
  AOI221_X1 vscale_core_DW_cmp_0_U449 ( .B1(vscale_core_DW_cmp_0n469), .B2(vscale_core_DW_cmp_0n594), .C1(pipeline_md_a[4]), .C2(vscale_core_DW_cmp_0n468), .A(vscale_core_DW_cmp_0n590), .ZN(
        vscale_core_DW_cmp_0n585) );
  NOR2_X1 vscale_core_DW_cmp_0_U450 ( .A1(vscale_core_DW_cmp_0n500), .A2(pipeline_md_b[5]), .ZN(vscale_core_DW_cmp_0n590) );
  OAI21_X1 vscale_core_DW_cmp_0_U451 ( .B1(pipeline_md_b[2]), .B2(vscale_core_DW_cmp_0n502), .A(vscale_core_DW_cmp_0n595), .ZN(vscale_core_DW_cmp_0n594) );
  AOI21_X1 vscale_core_DW_cmp_0_U452 ( .B1(vscale_core_DW_cmp_0n596), .B2(vscale_core_DW_cmp_0n469), .A(vscale_core_DW_cmp_0n587), .ZN(vscale_core_DW_cmp_0n584) );
  OAI21_X1 vscale_core_DW_cmp_0_U453 ( .B1(pipeline_md_b[6]), .B2(vscale_core_DW_cmp_0n503), .A(vscale_core_DW_cmp_0n593), .ZN(vscale_core_DW_cmp_0n587) );
  NAND2_X1 vscale_core_DW_cmp_0_U454 ( .A1(pipeline_md_a[7]), .A2(vscale_core_DW_cmp_0n467), .ZN(vscale_core_DW_cmp_0n593) );
  OAI21_X1 vscale_core_DW_cmp_0_U455 ( .B1(pipeline_md_a[3]), .B2(vscale_core_DW_cmp_0n470), .A(vscale_core_DW_cmp_0n598), .ZN(vscale_core_DW_cmp_0n597) );
  NAND3_X1 vscale_core_DW_cmp_0_U456 ( .A1(vscale_core_DW_cmp_0n595), .A2(vscale_core_DW_cmp_0n502), .A3(pipeline_md_b[2]), .ZN(vscale_core_DW_cmp_0n598) );
  NAND2_X1 vscale_core_DW_cmp_0_U457 ( .A1(pipeline_md_a[3]), .A2(vscale_core_DW_cmp_0n470), .ZN(vscale_core_DW_cmp_0n595) );
  AOI22_X1 vscale_core_DW_cmp_0_U458 ( .A1(pipeline_md_b[1]), .A2(vscale_core_DW_cmp_0n501), .B1(vscale_core_DW_cmp_0n599), .B2(pipeline_md_b[0]), .ZN(vscale_core_DW_cmp_0n596) );
  AOI21_X1 vscale_core_DW_cmp_0_U459 ( .B1(pipeline_md_a[1]), .B2(vscale_core_DW_cmp_0n471), .A(pipeline_md_a[0]), .ZN(vscale_core_DW_cmp_0n599) );
  OAI211_X1 vscale_core_DW_cmp_0_U460 ( .C1(pipeline_md_b[8]), .C2(vscale_core_DW_cmp_0n504), .A(vscale_core_DW_cmp_0n600), .B(vscale_core_DW_cmp_0n601), .ZN(vscale_core_DW_cmp_0n582) );
  NOR2_X1 vscale_core_DW_cmp_0_U461 ( .A1(vscale_core_DW_cmp_0n602), .A2(vscale_core_DW_cmp_0n603), .ZN(vscale_core_DW_cmp_0n601) );
  OAI21_X1 vscale_core_DW_cmp_0_U462 ( .B1(vscale_core_DW_cmp_0n602), .B2(vscale_core_DW_cmp_0n605), .A(vscale_core_DW_cmp_0n606), .ZN(vscale_core_DW_cmp_0n604) );
  OAI22_X1 vscale_core_DW_cmp_0_U463 ( .A1(vscale_core_DW_cmp_0n607), .A2(vscale_core_DW_cmp_0n608), .B1(vscale_core_DW_cmp_0n460), .B2(vscale_core_DW_cmp_0n607), .ZN(vscale_core_DW_cmp_0n606) );
  OAI21_X1 vscale_core_DW_cmp_0_U464 ( .B1(pipeline_md_a[13]), .B2(vscale_core_DW_cmp_0n462), .A(vscale_core_DW_cmp_0n609), .ZN(vscale_core_DW_cmp_0n608) );
  NAND3_X1 vscale_core_DW_cmp_0_U465 ( .A1(vscale_core_DW_cmp_0n610), .A2(vscale_core_DW_cmp_0n506), .A3(pipeline_md_b[12]), .ZN(vscale_core_DW_cmp_0n609) );
  OAI21_X1 vscale_core_DW_cmp_0_U466 ( .B1(pipeline_md_a[15]), .B2(vscale_core_DW_cmp_0n461), .A(vscale_core_DW_cmp_0n611), .ZN(vscale_core_DW_cmp_0n607) );
  NAND3_X1 vscale_core_DW_cmp_0_U467 ( .A1(vscale_core_DW_cmp_0n612), .A2(vscale_core_DW_cmp_0n507), .A3(pipeline_md_b[14]), .ZN(vscale_core_DW_cmp_0n611) );
  OAI22_X1 vscale_core_DW_cmp_0_U468 ( .A1(vscale_core_DW_cmp_0n613), .A2(vscale_core_DW_cmp_0n614), .B1(vscale_core_DW_cmp_0n463), .B2(vscale_core_DW_cmp_0n613), .ZN(vscale_core_DW_cmp_0n605) );
  OAI21_X1 vscale_core_DW_cmp_0_U469 ( .B1(pipeline_md_b[10]), .B2(vscale_core_DW_cmp_0n505), .A(vscale_core_DW_cmp_0n615), .ZN(vscale_core_DW_cmp_0n603) );
  OAI21_X1 vscale_core_DW_cmp_0_U470 ( .B1(pipeline_md_a[9]), .B2(vscale_core_DW_cmp_0n465), .A(vscale_core_DW_cmp_0n616), .ZN(vscale_core_DW_cmp_0n614) );
  NAND3_X1 vscale_core_DW_cmp_0_U471 ( .A1(vscale_core_DW_cmp_0n600), .A2(vscale_core_DW_cmp_0n504), .A3(pipeline_md_b[8]), .ZN(vscale_core_DW_cmp_0n616) );
  NAND2_X1 vscale_core_DW_cmp_0_U472 ( .A1(pipeline_md_a[9]), .A2(vscale_core_DW_cmp_0n465), .ZN(vscale_core_DW_cmp_0n600) );
  OAI21_X1 vscale_core_DW_cmp_0_U473 ( .B1(pipeline_md_a[11]), .B2(vscale_core_DW_cmp_0n464), .A(vscale_core_DW_cmp_0n617), .ZN(vscale_core_DW_cmp_0n613) );
  NAND3_X1 vscale_core_DW_cmp_0_U474 ( .A1(vscale_core_DW_cmp_0n615), .A2(vscale_core_DW_cmp_0n505), .A3(pipeline_md_b[10]), .ZN(vscale_core_DW_cmp_0n617) );
  NAND2_X1 vscale_core_DW_cmp_0_U475 ( .A1(pipeline_md_a[11]), .A2(vscale_core_DW_cmp_0n464), .ZN(vscale_core_DW_cmp_0n615) );
  OAI211_X1 vscale_core_DW_cmp_0_U476 ( .C1(pipeline_md_b[12]), .C2(vscale_core_DW_cmp_0n506), .A(vscale_core_DW_cmp_0n610), .B(vscale_core_DW_cmp_0n460), .ZN(vscale_core_DW_cmp_0n602) );
  OAI21_X1 vscale_core_DW_cmp_0_U477 ( .B1(pipeline_md_b[14]), .B2(vscale_core_DW_cmp_0n507), .A(vscale_core_DW_cmp_0n612), .ZN(vscale_core_DW_cmp_0n618) );
  NAND2_X1 vscale_core_DW_cmp_0_U478 ( .A1(pipeline_md_a[15]), .A2(vscale_core_DW_cmp_0n461), .ZN(vscale_core_DW_cmp_0n612) );
  NAND2_X1 vscale_core_DW_cmp_0_U479 ( .A1(pipeline_md_a[13]), .A2(vscale_core_DW_cmp_0n462), .ZN(vscale_core_DW_cmp_0n610) );
  NAND2_X1 vscale_core_DW_cmp_0_U480 ( .A1(pipeline_md_a[17]), .A2(vscale_core_DW_cmp_0n458), .ZN(vscale_core_DW_cmp_0n559) );
  OAI21_X1 vscale_core_DW_cmp_0_U481 ( .B1(vscale_core_DW_cmp_0n472), .B2(vscale_core_DW_cmp_0n619), .A(vscale_core_DW_cmp_0n620), .ZN(vscale_core_DW_cmp_0n531) );
  OAI22_X1 vscale_core_DW_cmp_0_U482 ( .A1(vscale_core_DW_cmp_0n621), .A2(vscale_core_DW_cmp_0n622), .B1(vscale_core_DW_cmp_0n473), .B2(vscale_core_DW_cmp_0n621), .ZN(vscale_core_DW_cmp_0n620) );
  OAI21_X1 vscale_core_DW_cmp_0_U483 ( .B1(vscale_core_DW_cmp_0n624), .B2(vscale_core_DW_cmp_0n625), .A(vscale_core_DW_cmp_0n626), .ZN(vscale_core_DW_cmp_0n622) );
  OAI22_X1 vscale_core_DW_cmp_0_U484 ( .A1(vscale_core_DW_cmp_0n627), .A2(vscale_core_DW_cmp_0n628), .B1(vscale_core_DW_cmp_0n494), .B2(vscale_core_DW_cmp_0n627), .ZN(vscale_core_DW_cmp_0n626) );
  OAI21_X1 vscale_core_DW_cmp_0_U485 ( .B1(pipeline_md_a[53]), .B2(vscale_core_DW_cmp_0n515), .A(vscale_core_DW_cmp_0n629), .ZN(vscale_core_DW_cmp_0n628) );
  NAND3_X1 vscale_core_DW_cmp_0_U486 ( .A1(vscale_core_DW_cmp_0n630), .A2(vscale_core_DW_cmp_0n493), .A3(pipeline_md_b[52]), .ZN(vscale_core_DW_cmp_0n629) );
  OAI21_X1 vscale_core_DW_cmp_0_U487 ( .B1(pipeline_md_a[55]), .B2(vscale_core_DW_cmp_0n514), .A(vscale_core_DW_cmp_0n631), .ZN(vscale_core_DW_cmp_0n627) );
  NAND3_X1 vscale_core_DW_cmp_0_U488 ( .A1(vscale_core_DW_cmp_0n632), .A2(vscale_core_DW_cmp_0n495), .A3(pipeline_md_b[54]), .ZN(vscale_core_DW_cmp_0n631) );
  OAI22_X1 vscale_core_DW_cmp_0_U489 ( .A1(vscale_core_DW_cmp_0n633), .A2(vscale_core_DW_cmp_0n634), .B1(vscale_core_DW_cmp_0n491), .B2(vscale_core_DW_cmp_0n633), .ZN(vscale_core_DW_cmp_0n625) );
  OAI21_X1 vscale_core_DW_cmp_0_U490 ( .B1(pipeline_md_a[49]), .B2(vscale_core_DW_cmp_0n517), .A(vscale_core_DW_cmp_0n636), .ZN(vscale_core_DW_cmp_0n634) );
  NAND3_X1 vscale_core_DW_cmp_0_U491 ( .A1(vscale_core_DW_cmp_0n637), .A2(vscale_core_DW_cmp_0n490), .A3(pipeline_md_b[48]), .ZN(vscale_core_DW_cmp_0n636) );
  OAI21_X1 vscale_core_DW_cmp_0_U492 ( .B1(pipeline_md_a[51]), .B2(vscale_core_DW_cmp_0n516), .A(vscale_core_DW_cmp_0n638), .ZN(vscale_core_DW_cmp_0n633) );
  NAND3_X1 vscale_core_DW_cmp_0_U493 ( .A1(vscale_core_DW_cmp_0n639), .A2(vscale_core_DW_cmp_0n492), .A3(pipeline_md_b[50]), .ZN(vscale_core_DW_cmp_0n638) );
  OAI22_X1 vscale_core_DW_cmp_0_U494 ( .A1(vscale_core_DW_cmp_0n640), .A2(vscale_core_DW_cmp_0n641), .B1(vscale_core_DW_cmp_0n474), .B2(vscale_core_DW_cmp_0n642), .ZN(vscale_core_DW_cmp_0n621) );
  OAI22_X1 vscale_core_DW_cmp_0_U495 ( .A1(vscale_core_DW_cmp_0n643), .A2(vscale_core_DW_cmp_0n644), .B1(vscale_core_DW_cmp_0n497), .B2(vscale_core_DW_cmp_0n643), .ZN(vscale_core_DW_cmp_0n642) );
  OAI21_X1 vscale_core_DW_cmp_0_U496 ( .B1(pipeline_md_a[57]), .B2(vscale_core_DW_cmp_0n513), .A(vscale_core_DW_cmp_0n646), .ZN(vscale_core_DW_cmp_0n644) );
  NAND3_X1 vscale_core_DW_cmp_0_U497 ( .A1(vscale_core_DW_cmp_0n647), .A2(vscale_core_DW_cmp_0n496), .A3(pipeline_md_b[56]), .ZN(vscale_core_DW_cmp_0n646) );
  OAI21_X1 vscale_core_DW_cmp_0_U498 ( .B1(pipeline_md_a[59]), .B2(vscale_core_DW_cmp_0n512), .A(vscale_core_DW_cmp_0n648), .ZN(vscale_core_DW_cmp_0n643) );
  NAND3_X1 vscale_core_DW_cmp_0_U499 ( .A1(vscale_core_DW_cmp_0n649), .A2(vscale_core_DW_cmp_0n498), .A3(pipeline_md_b[58]), .ZN(vscale_core_DW_cmp_0n648) );
  AOI221_X1 vscale_core_DW_cmp_0_U500 ( .B1(pipeline_md_b[62]), .B2(vscale_core_DW_cmp_0n530), .C1(pipeline_md_b[61]), .C2(vscale_core_DW_cmp_0n499), .A(vscale_core_DW_cmp_0n650), 
        .ZN(vscale_core_DW_cmp_0n640) );
  NOR3_X1 vscale_core_DW_cmp_0_U501 ( .A1(vscale_core_DW_cmp_0n511), .A2(pipeline_md_a[60]), .A3(vscale_core_DW_cmp_0n651), .ZN(vscale_core_DW_cmp_0n650) );
  OAI22_X1 vscale_core_DW_cmp_0_U502 ( .A1(vscale_core_DW_cmp_0n652), .A2(vscale_core_DW_cmp_0n653), .B1(vscale_core_DW_cmp_0n483), .B2(vscale_core_DW_cmp_0n652), .ZN(vscale_core_DW_cmp_0n619) );
  OAI211_X1 vscale_core_DW_cmp_0_U503 ( .C1(pipeline_md_b[40]), .C2(vscale_core_DW_cmp_0n484), .A(vscale_core_DW_cmp_0n654), .B(vscale_core_DW_cmp_0n655), .ZN(vscale_core_DW_cmp_0n537) );
  NOR2_X1 vscale_core_DW_cmp_0_U504 ( .A1(vscale_core_DW_cmp_0n656), .A2(vscale_core_DW_cmp_0n657), .ZN(vscale_core_DW_cmp_0n655) );
  OAI21_X1 vscale_core_DW_cmp_0_U505 ( .B1(vscale_core_DW_cmp_0n536), .B2(vscale_core_DW_cmp_0n658), .A(vscale_core_DW_cmp_0n659), .ZN(vscale_core_DW_cmp_0n653) );
  OAI22_X1 vscale_core_DW_cmp_0_U506 ( .A1(vscale_core_DW_cmp_0n660), .A2(vscale_core_DW_cmp_0n661), .B1(vscale_core_DW_cmp_0n481), .B2(vscale_core_DW_cmp_0n660), .ZN(vscale_core_DW_cmp_0n659) );
  OAI21_X1 vscale_core_DW_cmp_0_U507 ( .B1(pipeline_md_a[37]), .B2(vscale_core_DW_cmp_0n523), .A(vscale_core_DW_cmp_0n662), .ZN(vscale_core_DW_cmp_0n661) );
  NAND3_X1 vscale_core_DW_cmp_0_U508 ( .A1(vscale_core_DW_cmp_0n663), .A2(vscale_core_DW_cmp_0n480), .A3(pipeline_md_b[36]), .ZN(vscale_core_DW_cmp_0n662) );
  OAI21_X1 vscale_core_DW_cmp_0_U509 ( .B1(pipeline_md_a[39]), .B2(vscale_core_DW_cmp_0n522), .A(vscale_core_DW_cmp_0n664), .ZN(vscale_core_DW_cmp_0n660) );
  NAND3_X1 vscale_core_DW_cmp_0_U510 ( .A1(vscale_core_DW_cmp_0n665), .A2(vscale_core_DW_cmp_0n482), .A3(pipeline_md_b[38]), .ZN(vscale_core_DW_cmp_0n664) );
  OAI22_X1 vscale_core_DW_cmp_0_U511 ( .A1(vscale_core_DW_cmp_0n666), .A2(vscale_core_DW_cmp_0n667), .B1(vscale_core_DW_cmp_0n478), .B2(vscale_core_DW_cmp_0n666), .ZN(vscale_core_DW_cmp_0n658) );
  OAI21_X1 vscale_core_DW_cmp_0_U512 ( .B1(pipeline_md_b[34]), .B2(vscale_core_DW_cmp_0n479), .A(vscale_core_DW_cmp_0n668), .ZN(vscale_core_DW_cmp_0n535) );
  OAI21_X1 vscale_core_DW_cmp_0_U513 ( .B1(pipeline_md_a[33]), .B2(vscale_core_DW_cmp_0n525), .A(vscale_core_DW_cmp_0n669), .ZN(vscale_core_DW_cmp_0n667) );
  NAND3_X1 vscale_core_DW_cmp_0_U514 ( .A1(vscale_core_DW_cmp_0n538), .A2(vscale_core_DW_cmp_0n477), .A3(pipeline_md_b[32]), .ZN(vscale_core_DW_cmp_0n669) );
  NAND2_X1 vscale_core_DW_cmp_0_U515 ( .A1(pipeline_md_a[33]), .A2(vscale_core_DW_cmp_0n525), .ZN(vscale_core_DW_cmp_0n538) );
  OAI21_X1 vscale_core_DW_cmp_0_U516 ( .B1(pipeline_md_a[35]), .B2(vscale_core_DW_cmp_0n524), .A(vscale_core_DW_cmp_0n670), .ZN(vscale_core_DW_cmp_0n666) );
  NAND3_X1 vscale_core_DW_cmp_0_U517 ( .A1(vscale_core_DW_cmp_0n668), .A2(vscale_core_DW_cmp_0n479), .A3(pipeline_md_b[34]), .ZN(vscale_core_DW_cmp_0n670) );
  NAND2_X1 vscale_core_DW_cmp_0_U518 ( .A1(pipeline_md_a[35]), .A2(vscale_core_DW_cmp_0n524), .ZN(vscale_core_DW_cmp_0n668) );
  OAI211_X1 vscale_core_DW_cmp_0_U519 ( .C1(pipeline_md_b[36]), .C2(vscale_core_DW_cmp_0n480), .A(vscale_core_DW_cmp_0n663), .B(vscale_core_DW_cmp_0n481), .ZN(vscale_core_DW_cmp_0n536) );
  OAI21_X1 vscale_core_DW_cmp_0_U520 ( .B1(pipeline_md_b[38]), .B2(vscale_core_DW_cmp_0n482), .A(vscale_core_DW_cmp_0n665), .ZN(vscale_core_DW_cmp_0n671) );
  NAND2_X1 vscale_core_DW_cmp_0_U521 ( .A1(pipeline_md_a[39]), .A2(vscale_core_DW_cmp_0n522), .ZN(vscale_core_DW_cmp_0n665) );
  NAND2_X1 vscale_core_DW_cmp_0_U522 ( .A1(pipeline_md_a[37]), .A2(vscale_core_DW_cmp_0n523), .ZN(vscale_core_DW_cmp_0n663) );
  OAI21_X1 vscale_core_DW_cmp_0_U523 ( .B1(vscale_core_DW_cmp_0n656), .B2(vscale_core_DW_cmp_0n672), .A(vscale_core_DW_cmp_0n673), .ZN(vscale_core_DW_cmp_0n652) );
  OAI22_X1 vscale_core_DW_cmp_0_U524 ( .A1(vscale_core_DW_cmp_0n674), .A2(vscale_core_DW_cmp_0n675), .B1(vscale_core_DW_cmp_0n488), .B2(vscale_core_DW_cmp_0n674), .ZN(vscale_core_DW_cmp_0n673) );
  OAI21_X1 vscale_core_DW_cmp_0_U525 ( .B1(pipeline_md_a[45]), .B2(vscale_core_DW_cmp_0n519), .A(vscale_core_DW_cmp_0n676), .ZN(vscale_core_DW_cmp_0n675) );
  NAND3_X1 vscale_core_DW_cmp_0_U526 ( .A1(vscale_core_DW_cmp_0n677), .A2(vscale_core_DW_cmp_0n487), .A3(pipeline_md_b[44]), .ZN(vscale_core_DW_cmp_0n676) );
  OAI21_X1 vscale_core_DW_cmp_0_U527 ( .B1(pipeline_md_a[47]), .B2(vscale_core_DW_cmp_0n518), .A(vscale_core_DW_cmp_0n678), .ZN(vscale_core_DW_cmp_0n674) );
  NAND3_X1 vscale_core_DW_cmp_0_U528 ( .A1(vscale_core_DW_cmp_0n679), .A2(vscale_core_DW_cmp_0n489), .A3(pipeline_md_b[46]), .ZN(vscale_core_DW_cmp_0n678) );
  OAI22_X1 vscale_core_DW_cmp_0_U529 ( .A1(vscale_core_DW_cmp_0n680), .A2(vscale_core_DW_cmp_0n681), .B1(vscale_core_DW_cmp_0n485), .B2(vscale_core_DW_cmp_0n680), .ZN(vscale_core_DW_cmp_0n672) );
  OAI21_X1 vscale_core_DW_cmp_0_U530 ( .B1(pipeline_md_b[42]), .B2(vscale_core_DW_cmp_0n486), .A(vscale_core_DW_cmp_0n682), .ZN(vscale_core_DW_cmp_0n657) );
  OAI21_X1 vscale_core_DW_cmp_0_U531 ( .B1(pipeline_md_a[41]), .B2(vscale_core_DW_cmp_0n521), .A(vscale_core_DW_cmp_0n683), .ZN(vscale_core_DW_cmp_0n681) );
  NAND3_X1 vscale_core_DW_cmp_0_U532 ( .A1(vscale_core_DW_cmp_0n654), .A2(vscale_core_DW_cmp_0n484), .A3(pipeline_md_b[40]), .ZN(vscale_core_DW_cmp_0n683) );
  NAND2_X1 vscale_core_DW_cmp_0_U533 ( .A1(pipeline_md_a[41]), .A2(vscale_core_DW_cmp_0n521), .ZN(vscale_core_DW_cmp_0n654) );
  OAI21_X1 vscale_core_DW_cmp_0_U534 ( .B1(pipeline_md_a[43]), .B2(vscale_core_DW_cmp_0n520), .A(vscale_core_DW_cmp_0n684), .ZN(vscale_core_DW_cmp_0n680) );
  NAND3_X1 vscale_core_DW_cmp_0_U535 ( .A1(vscale_core_DW_cmp_0n682), .A2(vscale_core_DW_cmp_0n486), .A3(pipeline_md_b[42]), .ZN(vscale_core_DW_cmp_0n684) );
  NAND2_X1 vscale_core_DW_cmp_0_U536 ( .A1(pipeline_md_a[43]), .A2(vscale_core_DW_cmp_0n520), .ZN(vscale_core_DW_cmp_0n682) );
  OAI211_X1 vscale_core_DW_cmp_0_U537 ( .C1(pipeline_md_b[44]), .C2(vscale_core_DW_cmp_0n487), .A(vscale_core_DW_cmp_0n677), .B(vscale_core_DW_cmp_0n488), .ZN(vscale_core_DW_cmp_0n656) );
  OAI21_X1 vscale_core_DW_cmp_0_U538 ( .B1(pipeline_md_b[46]), .B2(vscale_core_DW_cmp_0n489), .A(vscale_core_DW_cmp_0n679), .ZN(vscale_core_DW_cmp_0n685) );
  NAND2_X1 vscale_core_DW_cmp_0_U539 ( .A1(pipeline_md_a[47]), .A2(vscale_core_DW_cmp_0n518), .ZN(vscale_core_DW_cmp_0n679) );
  NAND2_X1 vscale_core_DW_cmp_0_U540 ( .A1(pipeline_md_a[45]), .A2(vscale_core_DW_cmp_0n519), .ZN(vscale_core_DW_cmp_0n677) );
  NOR4_X1 vscale_core_DW_cmp_0_U541 ( .A1(vscale_core_DW_cmp_0n635), .A2(vscale_core_DW_cmp_0n623), .A3(vscale_core_DW_cmp_0n686), .A4(vscale_core_DW_cmp_0n624), .ZN(vscale_core_DW_cmp_0n539) );
  OAI211_X1 vscale_core_DW_cmp_0_U542 ( .C1(pipeline_md_b[52]), .C2(vscale_core_DW_cmp_0n493), .A(vscale_core_DW_cmp_0n630), .B(vscale_core_DW_cmp_0n494), .ZN(vscale_core_DW_cmp_0n624) );
  OAI21_X1 vscale_core_DW_cmp_0_U543 ( .B1(pipeline_md_b[54]), .B2(vscale_core_DW_cmp_0n495), .A(vscale_core_DW_cmp_0n632), .ZN(vscale_core_DW_cmp_0n687) );
  NAND2_X1 vscale_core_DW_cmp_0_U544 ( .A1(pipeline_md_a[55]), .A2(vscale_core_DW_cmp_0n514), .ZN(vscale_core_DW_cmp_0n632) );
  NAND2_X1 vscale_core_DW_cmp_0_U545 ( .A1(pipeline_md_a[53]), .A2(vscale_core_DW_cmp_0n515), .ZN(vscale_core_DW_cmp_0n630) );
  OAI21_X1 vscale_core_DW_cmp_0_U546 ( .B1(vscale_core_DW_cmp_0n490), .B2(pipeline_md_b[48]), .A(vscale_core_DW_cmp_0n637), .ZN(vscale_core_DW_cmp_0n686) );
  NAND2_X1 vscale_core_DW_cmp_0_U547 ( .A1(pipeline_md_a[49]), .A2(vscale_core_DW_cmp_0n517), .ZN(vscale_core_DW_cmp_0n637) );
  OAI211_X1 vscale_core_DW_cmp_0_U548 ( .C1(pipeline_md_b[56]), .C2(vscale_core_DW_cmp_0n496), .A(vscale_core_DW_cmp_0n647), .B(vscale_core_DW_cmp_0n688), .ZN(vscale_core_DW_cmp_0n623) );
  NOR2_X1 vscale_core_DW_cmp_0_U549 ( .A1(vscale_core_DW_cmp_0n474), .A2(vscale_core_DW_cmp_0n645), .ZN(vscale_core_DW_cmp_0n688) );
  OAI21_X1 vscale_core_DW_cmp_0_U550 ( .B1(pipeline_md_b[58]), .B2(vscale_core_DW_cmp_0n498), .A(vscale_core_DW_cmp_0n649), .ZN(vscale_core_DW_cmp_0n645) );
  NAND2_X1 vscale_core_DW_cmp_0_U551 ( .A1(pipeline_md_a[59]), .A2(vscale_core_DW_cmp_0n512), .ZN(vscale_core_DW_cmp_0n649) );
  AOI211_X1 vscale_core_DW_cmp_0_U552 ( .C1(vscale_core_DW_cmp_0n511), .C2(pipeline_md_a[60]), .A(vscale_core_DW_cmp_0n651), .B(vscale_core_DW_cmp_0n641), .ZN(vscale_core_DW_cmp_0n689) );
  OAI21_X1 vscale_core_DW_cmp_0_U553 ( .B1(pipeline_md_b[62]), .B2(vscale_core_DW_cmp_0n530), .A(vscale_core_DW_cmp_0n475), .ZN(vscale_core_DW_cmp_0n641) );
  NOR2_X1 vscale_core_DW_cmp_0_U554 ( .A1(vscale_core_DW_cmp_0n499), .A2(pipeline_md_b[61]), .ZN(vscale_core_DW_cmp_0n651) );
  NAND2_X1 vscale_core_DW_cmp_0_U555 ( .A1(pipeline_md_a[57]), .A2(vscale_core_DW_cmp_0n513), .ZN(vscale_core_DW_cmp_0n647) );
  OAI21_X1 vscale_core_DW_cmp_0_U556 ( .B1(pipeline_md_b[50]), .B2(vscale_core_DW_cmp_0n492), .A(vscale_core_DW_cmp_0n639), .ZN(vscale_core_DW_cmp_0n635) );
  NAND2_X1 vscale_core_DW_cmp_0_U557 ( .A1(pipeline_md_a[51]), .A2(vscale_core_DW_cmp_0n516), .ZN(vscale_core_DW_cmp_0n639) );
;
  vscale_core_DW01_sub_5 pipeline_md_sub_65 

  XOR2_X2 vscale_core_DW01_sub_5_U1 ( .A(vscale_core_DW01_sub_5n129), .B(vscale_core_DW01_sub_5n1), .Z(pipeline_md_N159) );
  HA_X1 vscale_core_DW01_sub_5_U2 ( .A(vscale_core_DW01_sub_5n130), .B(vscale_core_DW01_sub_5n2), .CO(vscale_core_DW01_sub_5n1), .S(pipeline_md_N158) );
  HA_X1 vscale_core_DW01_sub_5_U3 ( .A(vscale_core_DW01_sub_5n131), .B(vscale_core_DW01_sub_5n3), .CO(vscale_core_DW01_sub_5n2), .S(pipeline_md_N157) );
  HA_X1 vscale_core_DW01_sub_5_U4 ( .A(vscale_core_DW01_sub_5n132), .B(vscale_core_DW01_sub_5n4), .CO(vscale_core_DW01_sub_5n3), .S(pipeline_md_N156) );
  HA_X1 vscale_core_DW01_sub_5_U5 ( .A(vscale_core_DW01_sub_5n133), .B(vscale_core_DW01_sub_5n5), .CO(vscale_core_DW01_sub_5n4), .S(pipeline_md_N155) );
  HA_X1 vscale_core_DW01_sub_5_U6 ( .A(vscale_core_DW01_sub_5n134), .B(vscale_core_DW01_sub_5n6), .CO(vscale_core_DW01_sub_5n5), .S(pipeline_md_N154) );
  HA_X1 vscale_core_DW01_sub_5_U7 ( .A(vscale_core_DW01_sub_5n135), .B(vscale_core_DW01_sub_5n7), .CO(vscale_core_DW01_sub_5n6), .S(pipeline_md_N153) );
  HA_X1 vscale_core_DW01_sub_5_U8 ( .A(vscale_core_DW01_sub_5n136), .B(vscale_core_DW01_sub_5n8), .CO(vscale_core_DW01_sub_5n7), .S(pipeline_md_N152) );
  HA_X1 vscale_core_DW01_sub_5_U9 ( .A(vscale_core_DW01_sub_5n137), .B(vscale_core_DW01_sub_5n9), .CO(vscale_core_DW01_sub_5n8), .S(pipeline_md_N151) );
  HA_X1 vscale_core_DW01_sub_5_U10 ( .A(vscale_core_DW01_sub_5n138), .B(vscale_core_DW01_sub_5n10), .CO(vscale_core_DW01_sub_5n9), .S(pipeline_md_N150) );
  HA_X1 vscale_core_DW01_sub_5_U11 ( .A(vscale_core_DW01_sub_5n139), .B(vscale_core_DW01_sub_5n11), .CO(vscale_core_DW01_sub_5n10), .S(pipeline_md_N149) );
  HA_X1 vscale_core_DW01_sub_5_U12 ( .A(vscale_core_DW01_sub_5n140), .B(vscale_core_DW01_sub_5n12), .CO(vscale_core_DW01_sub_5n11), .S(pipeline_md_N148) );
  HA_X1 vscale_core_DW01_sub_5_U13 ( .A(vscale_core_DW01_sub_5n141), .B(vscale_core_DW01_sub_5n13), .CO(vscale_core_DW01_sub_5n12), .S(pipeline_md_N147) );
  HA_X1 vscale_core_DW01_sub_5_U14 ( .A(vscale_core_DW01_sub_5n142), .B(vscale_core_DW01_sub_5n14), .CO(vscale_core_DW01_sub_5n13), .S(pipeline_md_N146) );
  HA_X1 vscale_core_DW01_sub_5_U15 ( .A(vscale_core_DW01_sub_5n143), .B(vscale_core_DW01_sub_5n15), .CO(vscale_core_DW01_sub_5n14), .S(pipeline_md_N145) );
  HA_X1 vscale_core_DW01_sub_5_U16 ( .A(vscale_core_DW01_sub_5n144), .B(vscale_core_DW01_sub_5n16), .CO(vscale_core_DW01_sub_5n15), .S(pipeline_md_N144) );
  HA_X1 vscale_core_DW01_sub_5_U17 ( .A(vscale_core_DW01_sub_5n145), .B(vscale_core_DW01_sub_5n17), .CO(vscale_core_DW01_sub_5n16), .S(pipeline_md_N143) );
  HA_X1 vscale_core_DW01_sub_5_U18 ( .A(vscale_core_DW01_sub_5n146), .B(vscale_core_DW01_sub_5n18), .CO(vscale_core_DW01_sub_5n17), .S(pipeline_md_N142) );
  HA_X1 vscale_core_DW01_sub_5_U19 ( .A(vscale_core_DW01_sub_5n147), .B(vscale_core_DW01_sub_5n19), .CO(vscale_core_DW01_sub_5n18), .S(pipeline_md_N141) );
  HA_X1 vscale_core_DW01_sub_5_U20 ( .A(vscale_core_DW01_sub_5n148), .B(vscale_core_DW01_sub_5n346), .CO(vscale_core_DW01_sub_5n19), .S(pipeline_md_N140) );
  XNOR2_X2 vscale_core_DW01_sub_5_U22 ( .A(vscale_core_DW01_sub_5n22), .B(pipeline_md_result_muxed[43]), .ZN(pipeline_md_N139) );
  XNOR2_X2 vscale_core_DW01_sub_5_U25 ( .A(vscale_core_DW01_sub_5n25), .B(pipeline_md_result_muxed[42]), .ZN(pipeline_md_N138) );
  NAND2_X2 vscale_core_DW01_sub_5_U27 ( .A1(vscale_core_DW01_sub_5n33), .A2(vscale_core_DW01_sub_5n24), .ZN(vscale_core_DW01_sub_5n23) );
  XOR2_X2 vscale_core_DW01_sub_5_U29 ( .A(pipeline_md_result_muxed[41]), .B(vscale_core_DW01_sub_5n28), .Z(pipeline_md_N137) );
  NAND2_X2 vscale_core_DW01_sub_5_U31 ( .A1(vscale_core_DW01_sub_5n29), .A2(vscale_core_DW01_sub_5n27), .ZN(vscale_core_DW01_sub_5n26) );
  XOR2_X2 vscale_core_DW01_sub_5_U33 ( .A(pipeline_md_result_muxed[40]), .B(vscale_core_DW01_sub_5n30), .Z(pipeline_md_N136) );
  NAND2_X2 vscale_core_DW01_sub_5_U34 ( .A1(vscale_core_DW01_sub_5n31), .A2(vscale_core_DW01_sub_5n29), .ZN(vscale_core_DW01_sub_5n28) );
  XOR2_X2 vscale_core_DW01_sub_5_U36 ( .A(pipeline_md_result_muxed[39]), .B(vscale_core_DW01_sub_5n36), .Z(pipeline_md_N135) );
  NAND2_X2 vscale_core_DW01_sub_5_U41 ( .A1(vscale_core_DW01_sub_5n40), .A2(vscale_core_DW01_sub_5n35), .ZN(vscale_core_DW01_sub_5n34) );
  XNOR2_X2 vscale_core_DW01_sub_5_U43 ( .A(vscale_core_DW01_sub_5n38), .B(pipeline_md_result_muxed[38]), .ZN(pipeline_md_N134) );
  NAND2_X2 vscale_core_DW01_sub_5_U44 ( .A1(vscale_core_DW01_sub_5n38), .A2(vscale_core_DW01_sub_5n37), .ZN(vscale_core_DW01_sub_5n36) );
  XOR2_X2 vscale_core_DW01_sub_5_U46 ( .A(pipeline_md_result_muxed[37]), .B(vscale_core_DW01_sub_5n41), .Z(pipeline_md_N133) );
  XOR2_X2 vscale_core_DW01_sub_5_U50 ( .A(pipeline_md_result_muxed[36]), .B(vscale_core_DW01_sub_5n43), .Z(pipeline_md_N132) );
  NAND2_X2 vscale_core_DW01_sub_5_U51 ( .A1(vscale_core_DW01_sub_5n44), .A2(vscale_core_DW01_sub_5n42), .ZN(vscale_core_DW01_sub_5n41) );
  XOR2_X2 vscale_core_DW01_sub_5_U53 ( .A(pipeline_md_result_muxed[35]), .B(vscale_core_DW01_sub_5n47), .Z(pipeline_md_N131) );
  NAND2_X2 vscale_core_DW01_sub_5_U56 ( .A1(vscale_core_DW01_sub_5n51), .A2(vscale_core_DW01_sub_5n46), .ZN(vscale_core_DW01_sub_5n45) );
  XNOR2_X2 vscale_core_DW01_sub_5_U58 ( .A(vscale_core_DW01_sub_5n49), .B(pipeline_md_result_muxed[34]), .ZN(pipeline_md_N130) );
  NAND2_X2 vscale_core_DW01_sub_5_U59 ( .A1(vscale_core_DW01_sub_5n49), .A2(vscale_core_DW01_sub_5n48), .ZN(vscale_core_DW01_sub_5n47) );
  XNOR2_X2 vscale_core_DW01_sub_5_U61 ( .A(vscale_core_DW01_sub_5n52), .B(pipeline_md_result_muxed[33]), .ZN(pipeline_md_N129) );
  XOR2_X2 vscale_core_DW01_sub_5_U65 ( .A(pipeline_md_result_muxed[32]), .B(vscale_core_DW01_sub_5n53), .Z(pipeline_md_N128) );
  XNOR2_X2 vscale_core_DW01_sub_5_U67 ( .A(vscale_core_DW01_sub_5n59), .B(pipeline_md_result_muxed[31]), .ZN(pipeline_md_N127) );
  NAND2_X2 vscale_core_DW01_sub_5_U70 ( .A1(vscale_core_DW01_sub_5n74), .A2(vscale_core_DW01_sub_5n56), .ZN(vscale_core_DW01_sub_5n55) );
  NAND2_X2 vscale_core_DW01_sub_5_U72 ( .A1(vscale_core_DW01_sub_5n61), .A2(vscale_core_DW01_sub_5n58), .ZN(vscale_core_DW01_sub_5n57) );
  XOR2_X2 vscale_core_DW01_sub_5_U74 ( .A(pipeline_md_result_muxed[30]), .B(vscale_core_DW01_sub_5n60), .Z(pipeline_md_N126) );
  XNOR2_X2 vscale_core_DW01_sub_5_U76 ( .A(vscale_core_DW01_sub_5n62), .B(pipeline_md_result_muxed[29]), .ZN(pipeline_md_N125) );
  NAND2_X2 vscale_core_DW01_sub_5_U77 ( .A1(vscale_core_DW01_sub_5n63), .A2(vscale_core_DW01_sub_5n61), .ZN(vscale_core_DW01_sub_5n60) );
  XNOR2_X2 vscale_core_DW01_sub_5_U79 ( .A(vscale_core_DW01_sub_5n63), .B(pipeline_md_result_muxed[28]), .ZN(pipeline_md_N124) );
  XNOR2_X2 vscale_core_DW01_sub_5_U81 ( .A(vscale_core_DW01_sub_5n68), .B(pipeline_md_result_muxed[27]), .ZN(pipeline_md_N123) );
  NAND2_X2 vscale_core_DW01_sub_5_U83 ( .A1(vscale_core_DW01_sub_5n72), .A2(vscale_core_DW01_sub_5n65), .ZN(vscale_core_DW01_sub_5n64) );
  NAND2_X2 vscale_core_DW01_sub_5_U85 ( .A1(vscale_core_DW01_sub_5n70), .A2(vscale_core_DW01_sub_5n67), .ZN(vscale_core_DW01_sub_5n66) );
  XOR2_X2 vscale_core_DW01_sub_5_U87 ( .A(pipeline_md_result_muxed[26]), .B(vscale_core_DW01_sub_5n69), .Z(pipeline_md_N122) );
  XNOR2_X2 vscale_core_DW01_sub_5_U89 ( .A(vscale_core_DW01_sub_5n71), .B(pipeline_md_result_muxed[25]), .ZN(pipeline_md_N121) );
  NAND2_X2 vscale_core_DW01_sub_5_U90 ( .A1(vscale_core_DW01_sub_5n72), .A2(vscale_core_DW01_sub_5n70), .ZN(vscale_core_DW01_sub_5n69) );
  XNOR2_X2 vscale_core_DW01_sub_5_U92 ( .A(vscale_core_DW01_sub_5n72), .B(pipeline_md_result_muxed[24]), .ZN(pipeline_md_N120) );
  XNOR2_X2 vscale_core_DW01_sub_5_U94 ( .A(vscale_core_DW01_sub_5n77), .B(pipeline_md_result_muxed[23]), .ZN(pipeline_md_N119) );
  NAND2_X2 vscale_core_DW01_sub_5_U96 ( .A1(vscale_core_DW01_sub_5n91), .A2(vscale_core_DW01_sub_5n74), .ZN(vscale_core_DW01_sub_5n73) );
  NAND2_X2 vscale_core_DW01_sub_5_U98 ( .A1(vscale_core_DW01_sub_5n79), .A2(vscale_core_DW01_sub_5n76), .ZN(vscale_core_DW01_sub_5n75) );
  XOR2_X2 vscale_core_DW01_sub_5_U100 ( .A(pipeline_md_result_muxed[22]), .B(vscale_core_DW01_sub_5n78), .Z(pipeline_md_N118) );
  XNOR2_X2 vscale_core_DW01_sub_5_U102 ( .A(vscale_core_DW01_sub_5n80), .B(pipeline_md_result_muxed[21]), .ZN(pipeline_md_N117) );
  NAND2_X2 vscale_core_DW01_sub_5_U103 ( .A1(vscale_core_DW01_sub_5n81), .A2(vscale_core_DW01_sub_5n79), .ZN(vscale_core_DW01_sub_5n78) );
  XNOR2_X2 vscale_core_DW01_sub_5_U105 ( .A(vscale_core_DW01_sub_5n81), .B(pipeline_md_result_muxed[20]), .ZN(pipeline_md_N116) );
  XNOR2_X2 vscale_core_DW01_sub_5_U107 ( .A(vscale_core_DW01_sub_5n86), .B(pipeline_md_result_muxed[19]), .ZN(pipeline_md_N115) );
  NAND2_X2 vscale_core_DW01_sub_5_U109 ( .A1(vscale_core_DW01_sub_5n91), .A2(vscale_core_DW01_sub_5n83), .ZN(vscale_core_DW01_sub_5n82) );
  NAND2_X2 vscale_core_DW01_sub_5_U111 ( .A1(vscale_core_DW01_sub_5n88), .A2(vscale_core_DW01_sub_5n85), .ZN(vscale_core_DW01_sub_5n84) );
  XOR2_X2 vscale_core_DW01_sub_5_U113 ( .A(pipeline_md_result_muxed[18]), .B(vscale_core_DW01_sub_5n87), .Z(pipeline_md_N114) );
  XOR2_X2 vscale_core_DW01_sub_5_U115 ( .A(pipeline_md_result_muxed[17]), .B(vscale_core_DW01_sub_5n89), .Z(pipeline_md_N113) );
  NAND2_X2 vscale_core_DW01_sub_5_U116 ( .A1(vscale_core_DW01_sub_5n91), .A2(vscale_core_DW01_sub_5n88), .ZN(vscale_core_DW01_sub_5n87) );
  XNOR2_X2 vscale_core_DW01_sub_5_U118 ( .A(vscale_core_DW01_sub_5n91), .B(pipeline_md_result_muxed[16]), .ZN(pipeline_md_N112) );
  NAND2_X2 vscale_core_DW01_sub_5_U119 ( .A1(vscale_core_DW01_sub_5n91), .A2(vscale_core_DW01_sub_5n90), .ZN(vscale_core_DW01_sub_5n89) );
  XOR2_X2 vscale_core_DW01_sub_5_U121 ( .A(pipeline_md_result_muxed[15]), .B(vscale_core_DW01_sub_5n96), .Z(pipeline_md_N111) );
  NAND2_X2 vscale_core_DW01_sub_5_U123 ( .A1(vscale_core_DW01_sub_5n93), .A2(vscale_core_DW01_sub_5n114), .ZN(vscale_core_DW01_sub_5n92) );
  NAND2_X2 vscale_core_DW01_sub_5_U125 ( .A1(vscale_core_DW01_sub_5n100), .A2(vscale_core_DW01_sub_5n95), .ZN(vscale_core_DW01_sub_5n94) );
  XNOR2_X2 vscale_core_DW01_sub_5_U127 ( .A(vscale_core_DW01_sub_5n98), .B(pipeline_md_result_muxed[14]), .ZN(pipeline_md_N110) );
  NAND2_X2 vscale_core_DW01_sub_5_U128 ( .A1(vscale_core_DW01_sub_5n98), .A2(vscale_core_DW01_sub_5n97), .ZN(vscale_core_DW01_sub_5n96) );
  XOR2_X2 vscale_core_DW01_sub_5_U130 ( .A(pipeline_md_result_muxed[13]), .B(vscale_core_DW01_sub_5n101), .Z(pipeline_md_N109) );
  XOR2_X2 vscale_core_DW01_sub_5_U134 ( .A(pipeline_md_result_muxed[12]), .B(vscale_core_DW01_sub_5n103), .Z(pipeline_md_N108) );
  NAND2_X2 vscale_core_DW01_sub_5_U135 ( .A1(vscale_core_DW01_sub_5n104), .A2(vscale_core_DW01_sub_5n102), .ZN(vscale_core_DW01_sub_5n101) );
  XOR2_X2 vscale_core_DW01_sub_5_U137 ( .A(pipeline_md_result_muxed[11]), .B(vscale_core_DW01_sub_5n107), .Z(pipeline_md_N107) );
  NAND2_X2 vscale_core_DW01_sub_5_U140 ( .A1(vscale_core_DW01_sub_5n111), .A2(vscale_core_DW01_sub_5n106), .ZN(vscale_core_DW01_sub_5n105) );
  XNOR2_X2 vscale_core_DW01_sub_5_U142 ( .A(vscale_core_DW01_sub_5n109), .B(pipeline_md_result_muxed[10]), .ZN(pipeline_md_N106) );
  NAND2_X2 vscale_core_DW01_sub_5_U143 ( .A1(vscale_core_DW01_sub_5n109), .A2(vscale_core_DW01_sub_5n108), .ZN(vscale_core_DW01_sub_5n107) );
  XNOR2_X2 vscale_core_DW01_sub_5_U145 ( .A(vscale_core_DW01_sub_5n112), .B(pipeline_md_result_muxed[9]), .ZN(pipeline_md_N105) );
  XOR2_X2 vscale_core_DW01_sub_5_U149 ( .A(pipeline_md_result_muxed[8]), .B(vscale_core_DW01_sub_5n113), .Z(pipeline_md_N104) );
  XNOR2_X2 vscale_core_DW01_sub_5_U151 ( .A(vscale_core_DW01_sub_5n117), .B(pipeline_md_result_muxed[7]), .ZN(pipeline_md_N103) );
  NAND2_X2 vscale_core_DW01_sub_5_U154 ( .A1(vscale_core_DW01_sub_5n119), .A2(vscale_core_DW01_sub_5n116), .ZN(vscale_core_DW01_sub_5n115) );
  XOR2_X2 vscale_core_DW01_sub_5_U156 ( .A(pipeline_md_result_muxed[6]), .B(vscale_core_DW01_sub_5n118), .Z(pipeline_md_N102) );
  XOR2_X2 vscale_core_DW01_sub_5_U158 ( .A(pipeline_md_result_muxed[5]), .B(vscale_core_DW01_sub_5n120), .Z(pipeline_md_N101) );
  NAND2_X2 vscale_core_DW01_sub_5_U159 ( .A1(vscale_core_DW01_sub_5n122), .A2(vscale_core_DW01_sub_5n119), .ZN(vscale_core_DW01_sub_5n118) );
  XNOR2_X2 vscale_core_DW01_sub_5_U161 ( .A(vscale_core_DW01_sub_5n122), .B(pipeline_md_result_muxed[4]), .ZN(pipeline_md_N100) );
  NAND2_X2 vscale_core_DW01_sub_5_U162 ( .A1(vscale_core_DW01_sub_5n122), .A2(vscale_core_DW01_sub_5n121), .ZN(vscale_core_DW01_sub_5n120) );
  XNOR2_X2 vscale_core_DW01_sub_5_U164 ( .A(vscale_core_DW01_sub_5n125), .B(pipeline_md_result_muxed[3]), .ZN(pipeline_md_N99) );
  NAND2_X2 vscale_core_DW01_sub_5_U166 ( .A1(vscale_core_DW01_sub_5n124), .A2(vscale_core_DW01_sub_5n127), .ZN(vscale_core_DW01_sub_5n123) );
  XOR2_X2 vscale_core_DW01_sub_5_U168 ( .A(pipeline_md_result_muxed[2]), .B(vscale_core_DW01_sub_5n126), .Z(pipeline_md_N98) );
  XOR2_X2 vscale_core_DW01_sub_5_U170 ( .A(pipeline_md_result_muxed[0]), .B(pipeline_md_result_muxed[1]), .Z(pipeline_md_N97) );
  AND2_X4 vscale_core_DW01_sub_5_U196 ( .A1(vscale_core_DW01_sub_5n54), .A2(vscale_core_DW01_sub_5n21), .ZN(vscale_core_DW01_sub_5n346) );
  NOR2_X2 vscale_core_DW01_sub_5_U197 ( .A1(vscale_core_DW01_sub_5n55), .A2(vscale_core_DW01_sub_5n92), .ZN(vscale_core_DW01_sub_5n54) );
  NOR2_X2 vscale_core_DW01_sub_5_U198 ( .A1(vscale_core_DW01_sub_5n66), .A2(vscale_core_DW01_sub_5n57), .ZN(vscale_core_DW01_sub_5n56) );
  NOR2_X2 vscale_core_DW01_sub_5_U199 ( .A1(vscale_core_DW01_sub_5n53), .A2(vscale_core_DW01_sub_5n45), .ZN(vscale_core_DW01_sub_5n44) );
  NOR2_X2 vscale_core_DW01_sub_5_U200 ( .A1(vscale_core_DW01_sub_5n53), .A2(vscale_core_DW01_sub_5n32), .ZN(vscale_core_DW01_sub_5n31) );
  NOR2_X2 vscale_core_DW01_sub_5_U201 ( .A1(vscale_core_DW01_sub_5n43), .A2(vscale_core_DW01_sub_5n39), .ZN(vscale_core_DW01_sub_5n38) );
  NOR2_X2 vscale_core_DW01_sub_5_U202 ( .A1(vscale_core_DW01_sub_5n53), .A2(vscale_core_DW01_sub_5n50), .ZN(vscale_core_DW01_sub_5n49) );
  NOR2_X2 vscale_core_DW01_sub_5_U203 ( .A1(vscale_core_DW01_sub_5n113), .A2(vscale_core_DW01_sub_5n105), .ZN(vscale_core_DW01_sub_5n104) );
  NOR2_X2 vscale_core_DW01_sub_5_U204 ( .A1(vscale_core_DW01_sub_5n103), .A2(vscale_core_DW01_sub_5n99), .ZN(vscale_core_DW01_sub_5n98) );
  NOR2_X2 vscale_core_DW01_sub_5_U205 ( .A1(vscale_core_DW01_sub_5n113), .A2(vscale_core_DW01_sub_5n110), .ZN(vscale_core_DW01_sub_5n109) );
  NOR2_X2 vscale_core_DW01_sub_5_U206 ( .A1(pipeline_md_result_muxed[34]), .A2(pipeline_md_result_muxed[35]), .ZN(vscale_core_DW01_sub_5n46) );
  NOR2_X2 vscale_core_DW01_sub_5_U207 ( .A1(vscale_core_DW01_sub_5n26), .A2(pipeline_md_result_muxed[42]), .ZN(vscale_core_DW01_sub_5n24) );
  NOR2_X2 vscale_core_DW01_sub_5_U208 ( .A1(vscale_core_DW01_sub_5n105), .A2(vscale_core_DW01_sub_5n94), .ZN(vscale_core_DW01_sub_5n93) );
  NOR2_X2 vscale_core_DW01_sub_5_U209 ( .A1(pipeline_md_result_muxed[14]), .A2(pipeline_md_result_muxed[15]), .ZN(vscale_core_DW01_sub_5n95) );
  NOR2_X2 vscale_core_DW01_sub_5_U210 ( .A1(pipeline_md_result_muxed[2]), .A2(pipeline_md_result_muxed[3]), .ZN(vscale_core_DW01_sub_5n124) );
  NOR2_X2 vscale_core_DW01_sub_5_U211 ( .A1(pipeline_md_result_muxed[32]), .A2(pipeline_md_result_muxed[33]), .ZN(vscale_core_DW01_sub_5n51) );
  NOR2_X2 vscale_core_DW01_sub_5_U212 ( .A1(pipeline_md_result_muxed[36]), .A2(pipeline_md_result_muxed[37]), .ZN(vscale_core_DW01_sub_5n40) );
  NOR2_X2 vscale_core_DW01_sub_5_U213 ( .A1(pipeline_md_result_muxed[8]), .A2(pipeline_md_result_muxed[9]), .ZN(vscale_core_DW01_sub_5n111) );
  NOR2_X2 vscale_core_DW01_sub_5_U214 ( .A1(pipeline_md_result_muxed[12]), .A2(pipeline_md_result_muxed[13]), .ZN(vscale_core_DW01_sub_5n100) );
  NOR2_X2 vscale_core_DW01_sub_5_U215 ( .A1(vscale_core_DW01_sub_5n45), .A2(vscale_core_DW01_sub_5n34), .ZN(vscale_core_DW01_sub_5n33) );
  NOR2_X2 vscale_core_DW01_sub_5_U216 ( .A1(pipeline_md_result_muxed[38]), .A2(pipeline_md_result_muxed[39]), .ZN(vscale_core_DW01_sub_5n35) );
  NOR2_X2 vscale_core_DW01_sub_5_U217 ( .A1(pipeline_md_result_muxed[1]), .A2(pipeline_md_result_muxed[0]), .ZN(vscale_core_DW01_sub_5n127) );
  NOR2_X2 vscale_core_DW01_sub_5_U218 ( .A1(vscale_core_DW01_sub_5n115), .A2(vscale_core_DW01_sub_5n123), .ZN(vscale_core_DW01_sub_5n114) );
  NOR2_X2 vscale_core_DW01_sub_5_U219 ( .A1(pipeline_md_result_muxed[6]), .A2(pipeline_md_result_muxed[7]), .ZN(vscale_core_DW01_sub_5n116) );
  NOR2_X2 vscale_core_DW01_sub_5_U220 ( .A1(pipeline_md_result_muxed[24]), .A2(pipeline_md_result_muxed[25]), .ZN(vscale_core_DW01_sub_5n70) );
  NOR2_X2 vscale_core_DW01_sub_5_U221 ( .A1(pipeline_md_result_muxed[28]), .A2(pipeline_md_result_muxed[29]), .ZN(vscale_core_DW01_sub_5n61) );
  NOR2_X2 vscale_core_DW01_sub_5_U222 ( .A1(pipeline_md_result_muxed[20]), .A2(pipeline_md_result_muxed[21]), .ZN(vscale_core_DW01_sub_5n79) );
  NOR2_X2 vscale_core_DW01_sub_5_U223 ( .A1(pipeline_md_result_muxed[4]), .A2(pipeline_md_result_muxed[5]), .ZN(vscale_core_DW01_sub_5n119) );
  NOR2_X2 vscale_core_DW01_sub_5_U224 ( .A1(pipeline_md_result_muxed[16]), .A2(pipeline_md_result_muxed[17]), .ZN(vscale_core_DW01_sub_5n88) );
  NOR2_X2 vscale_core_DW01_sub_5_U225 ( .A1(vscale_core_DW01_sub_5n84), .A2(vscale_core_DW01_sub_5n75), .ZN(vscale_core_DW01_sub_5n74) );
  NOR2_X2 vscale_core_DW01_sub_5_U226 ( .A1(pipeline_md_result_muxed[22]), .A2(pipeline_md_result_muxed[23]), .ZN(vscale_core_DW01_sub_5n76) );
  NOR2_X2 vscale_core_DW01_sub_5_U227 ( .A1(pipeline_md_result_muxed[30]), .A2(pipeline_md_result_muxed[31]), .ZN(vscale_core_DW01_sub_5n58) );
  NOR2_X2 vscale_core_DW01_sub_5_U228 ( .A1(pipeline_md_result_muxed[26]), .A2(pipeline_md_result_muxed[27]), .ZN(vscale_core_DW01_sub_5n67) );
  NOR2_X2 vscale_core_DW01_sub_5_U229 ( .A1(pipeline_md_result_muxed[18]), .A2(pipeline_md_result_muxed[19]), .ZN(vscale_core_DW01_sub_5n85) );
  NOR2_X2 vscale_core_DW01_sub_5_U230 ( .A1(pipeline_md_result_muxed[10]), .A2(pipeline_md_result_muxed[11]), .ZN(vscale_core_DW01_sub_5n106) );
  NOR2_X2 vscale_core_DW01_sub_5_U231 ( .A1(vscale_core_DW01_sub_5n23), .A2(pipeline_md_result_muxed[43]), .ZN(vscale_core_DW01_sub_5n21) );
  NOR2_X2 vscale_core_DW01_sub_5_U232 ( .A1(vscale_core_DW01_sub_5n30), .A2(vscale_core_DW01_sub_5n26), .ZN(vscale_core_DW01_sub_5n25) );
  NOR2_X2 vscale_core_DW01_sub_5_U233 ( .A1(vscale_core_DW01_sub_5n64), .A2(pipeline_md_result_muxed[28]), .ZN(vscale_core_DW01_sub_5n62) );
  NOR2_X2 vscale_core_DW01_sub_5_U234 ( .A1(vscale_core_DW01_sub_5n60), .A2(pipeline_md_result_muxed[30]), .ZN(vscale_core_DW01_sub_5n59) );
  NOR2_X2 vscale_core_DW01_sub_5_U235 ( .A1(vscale_core_DW01_sub_5n53), .A2(vscale_core_DW01_sub_5n23), .ZN(vscale_core_DW01_sub_5n22) );
  NOR2_X2 vscale_core_DW01_sub_5_U236 ( .A1(vscale_core_DW01_sub_5n53), .A2(pipeline_md_result_muxed[32]), .ZN(vscale_core_DW01_sub_5n52) );
  NOR2_X2 vscale_core_DW01_sub_5_U237 ( .A1(vscale_core_DW01_sub_5n73), .A2(pipeline_md_result_muxed[24]), .ZN(vscale_core_DW01_sub_5n71) );
  NOR2_X2 vscale_core_DW01_sub_5_U238 ( .A1(vscale_core_DW01_sub_5n82), .A2(pipeline_md_result_muxed[20]), .ZN(vscale_core_DW01_sub_5n80) );
  NOR2_X2 vscale_core_DW01_sub_5_U239 ( .A1(vscale_core_DW01_sub_5n69), .A2(pipeline_md_result_muxed[26]), .ZN(vscale_core_DW01_sub_5n68) );
  NOR2_X2 vscale_core_DW01_sub_5_U240 ( .A1(vscale_core_DW01_sub_5n78), .A2(pipeline_md_result_muxed[22]), .ZN(vscale_core_DW01_sub_5n77) );
  NOR2_X2 vscale_core_DW01_sub_5_U241 ( .A1(vscale_core_DW01_sub_5n87), .A2(pipeline_md_result_muxed[18]), .ZN(vscale_core_DW01_sub_5n86) );
  NOR2_X2 vscale_core_DW01_sub_5_U242 ( .A1(vscale_core_DW01_sub_5n113), .A2(pipeline_md_result_muxed[8]), .ZN(vscale_core_DW01_sub_5n112) );
  NOR2_X2 vscale_core_DW01_sub_5_U243 ( .A1(vscale_core_DW01_sub_5n118), .A2(pipeline_md_result_muxed[6]), .ZN(vscale_core_DW01_sub_5n117) );
  NOR2_X2 vscale_core_DW01_sub_5_U244 ( .A1(vscale_core_DW01_sub_5n126), .A2(pipeline_md_result_muxed[2]), .ZN(vscale_core_DW01_sub_5n125) );
  BUF_X4 vscale_core_DW01_sub_5_U245 ( .A(pipeline_md_result_muxed[0]), .Z(pipeline_md_N96) );
  INV_X4 vscale_core_DW01_sub_5_U246 ( .A(vscale_core_DW01_sub_5n100), .ZN(vscale_core_DW01_sub_5n99) );
  INV_X4 vscale_core_DW01_sub_5_U247 ( .A(pipeline_md_result_muxed[14]), .ZN(vscale_core_DW01_sub_5n97) );
  INV_X4 vscale_core_DW01_sub_5_U248 ( .A(vscale_core_DW01_sub_5n92), .ZN(vscale_core_DW01_sub_5n91) );
  INV_X4 vscale_core_DW01_sub_5_U249 ( .A(pipeline_md_result_muxed[16]), .ZN(vscale_core_DW01_sub_5n90) );
  INV_X4 vscale_core_DW01_sub_5_U250 ( .A(vscale_core_DW01_sub_5n84), .ZN(vscale_core_DW01_sub_5n83) );
  INV_X4 vscale_core_DW01_sub_5_U251 ( .A(vscale_core_DW01_sub_5n82), .ZN(vscale_core_DW01_sub_5n81) );
  INV_X4 vscale_core_DW01_sub_5_U252 ( .A(vscale_core_DW01_sub_5n73), .ZN(vscale_core_DW01_sub_5n72) );
  INV_X4 vscale_core_DW01_sub_5_U253 ( .A(vscale_core_DW01_sub_5n66), .ZN(vscale_core_DW01_sub_5n65) );
  INV_X4 vscale_core_DW01_sub_5_U254 ( .A(vscale_core_DW01_sub_5n64), .ZN(vscale_core_DW01_sub_5n63) );
  INV_X4 vscale_core_DW01_sub_5_U255 ( .A(vscale_core_DW01_sub_5n54), .ZN(vscale_core_DW01_sub_5n53) );
  INV_X4 vscale_core_DW01_sub_5_U256 ( .A(vscale_core_DW01_sub_5n51), .ZN(vscale_core_DW01_sub_5n50) );
  INV_X4 vscale_core_DW01_sub_5_U257 ( .A(pipeline_md_result_muxed[34]), .ZN(vscale_core_DW01_sub_5n48) );
  INV_X4 vscale_core_DW01_sub_5_U258 ( .A(vscale_core_DW01_sub_5n44), .ZN(vscale_core_DW01_sub_5n43) );
  INV_X4 vscale_core_DW01_sub_5_U259 ( .A(pipeline_md_result_muxed[36]), .ZN(vscale_core_DW01_sub_5n42) );
  INV_X4 vscale_core_DW01_sub_5_U260 ( .A(vscale_core_DW01_sub_5n40), .ZN(vscale_core_DW01_sub_5n39) );
  INV_X4 vscale_core_DW01_sub_5_U261 ( .A(pipeline_md_result_muxed[38]), .ZN(vscale_core_DW01_sub_5n37) );
  INV_X4 vscale_core_DW01_sub_5_U262 ( .A(vscale_core_DW01_sub_5n33), .ZN(vscale_core_DW01_sub_5n32) );
  INV_X4 vscale_core_DW01_sub_5_U263 ( .A(vscale_core_DW01_sub_5n31), .ZN(vscale_core_DW01_sub_5n30) );
  INV_X4 vscale_core_DW01_sub_5_U264 ( .A(pipeline_md_result_muxed[40]), .ZN(vscale_core_DW01_sub_5n29) );
  INV_X4 vscale_core_DW01_sub_5_U265 ( .A(pipeline_md_result_muxed[41]), .ZN(vscale_core_DW01_sub_5n27) );
  INV_X4 vscale_core_DW01_sub_5_U266 ( .A(pipeline_md_result_muxed[44]), .ZN(vscale_core_DW01_sub_5n148) );
  INV_X4 vscale_core_DW01_sub_5_U267 ( .A(pipeline_md_result_muxed[45]), .ZN(vscale_core_DW01_sub_5n147) );
  INV_X4 vscale_core_DW01_sub_5_U268 ( .A(pipeline_md_result_muxed[46]), .ZN(vscale_core_DW01_sub_5n146) );
  INV_X4 vscale_core_DW01_sub_5_U269 ( .A(pipeline_md_result_muxed[47]), .ZN(vscale_core_DW01_sub_5n145) );
  INV_X4 vscale_core_DW01_sub_5_U270 ( .A(pipeline_md_result_muxed[48]), .ZN(vscale_core_DW01_sub_5n144) );
  INV_X4 vscale_core_DW01_sub_5_U271 ( .A(pipeline_md_result_muxed[49]), .ZN(vscale_core_DW01_sub_5n143) );
  INV_X4 vscale_core_DW01_sub_5_U272 ( .A(pipeline_md_result_muxed[50]), .ZN(vscale_core_DW01_sub_5n142) );
  INV_X4 vscale_core_DW01_sub_5_U273 ( .A(pipeline_md_result_muxed[51]), .ZN(vscale_core_DW01_sub_5n141) );
  INV_X4 vscale_core_DW01_sub_5_U274 ( .A(pipeline_md_result_muxed[52]), .ZN(vscale_core_DW01_sub_5n140) );
  INV_X4 vscale_core_DW01_sub_5_U275 ( .A(pipeline_md_result_muxed[53]), .ZN(vscale_core_DW01_sub_5n139) );
  INV_X4 vscale_core_DW01_sub_5_U276 ( .A(pipeline_md_result_muxed[54]), .ZN(vscale_core_DW01_sub_5n138) );
  INV_X4 vscale_core_DW01_sub_5_U277 ( .A(pipeline_md_result_muxed[55]), .ZN(vscale_core_DW01_sub_5n137) );
  INV_X4 vscale_core_DW01_sub_5_U278 ( .A(pipeline_md_result_muxed[56]), .ZN(vscale_core_DW01_sub_5n136) );
  INV_X4 vscale_core_DW01_sub_5_U279 ( .A(pipeline_md_result_muxed[57]), .ZN(vscale_core_DW01_sub_5n135) );
  INV_X4 vscale_core_DW01_sub_5_U280 ( .A(pipeline_md_result_muxed[58]), .ZN(vscale_core_DW01_sub_5n134) );
  INV_X4 vscale_core_DW01_sub_5_U281 ( .A(pipeline_md_result_muxed[59]), .ZN(vscale_core_DW01_sub_5n133) );
  INV_X4 vscale_core_DW01_sub_5_U282 ( .A(pipeline_md_result_muxed[60]), .ZN(vscale_core_DW01_sub_5n132) );
  INV_X4 vscale_core_DW01_sub_5_U283 ( .A(pipeline_md_result_muxed[61]), .ZN(vscale_core_DW01_sub_5n131) );
  INV_X4 vscale_core_DW01_sub_5_U284 ( .A(pipeline_md_result_muxed[62]), .ZN(vscale_core_DW01_sub_5n130) );
  INV_X4 vscale_core_DW01_sub_5_U285 ( .A(pipeline_md_result_muxed[63]), .ZN(vscale_core_DW01_sub_5n129) );
  INV_X4 vscale_core_DW01_sub_5_U286 ( .A(vscale_core_DW01_sub_5n127), .ZN(vscale_core_DW01_sub_5n126) );
  INV_X4 vscale_core_DW01_sub_5_U287 ( .A(vscale_core_DW01_sub_5n123), .ZN(vscale_core_DW01_sub_5n122) );
  INV_X4 vscale_core_DW01_sub_5_U288 ( .A(pipeline_md_result_muxed[4]), .ZN(vscale_core_DW01_sub_5n121) );
  INV_X4 vscale_core_DW01_sub_5_U289 ( .A(vscale_core_DW01_sub_5n114), .ZN(vscale_core_DW01_sub_5n113) );
  INV_X4 vscale_core_DW01_sub_5_U290 ( .A(vscale_core_DW01_sub_5n111), .ZN(vscale_core_DW01_sub_5n110) );
  INV_X4 vscale_core_DW01_sub_5_U291 ( .A(pipeline_md_result_muxed[10]), .ZN(vscale_core_DW01_sub_5n108) );
  INV_X4 vscale_core_DW01_sub_5_U292 ( .A(vscale_core_DW01_sub_5n104), .ZN(vscale_core_DW01_sub_5n103) );
  INV_X4 vscale_core_DW01_sub_5_U293 ( .A(pipeline_md_result_muxed[12]), .ZN(vscale_core_DW01_sub_5n102) );
;
  vscale_core_DW01_sub_6 pipeline_md_sub_109 

  XNOR2_X2 vscale_core_DW01_sub_6_U1 ( .A(vscale_core_DW01_sub_6n54), .B(n10233), .ZN(pipeline_md_N314) );
  FA_X1 vscale_core_DW01_sub_6_U2 ( .A(vscale_core_DW01_sub_6n400), .B(pipeline_md_a[62]), .CI(vscale_core_DW01_sub_6n55), .CO(vscale_core_DW01_sub_6n54), .S(pipeline_md_N313) );
  FA_X1 vscale_core_DW01_sub_6_U3 ( .A(vscale_core_DW01_sub_6n401), .B(pipeline_md_a[61]), .CI(vscale_core_DW01_sub_6n56), .CO(vscale_core_DW01_sub_6n55), .S(pipeline_md_N312) );
  FA_X1 vscale_core_DW01_sub_6_U4 ( .A(vscale_core_DW01_sub_6n402), .B(pipeline_md_a[60]), .CI(vscale_core_DW01_sub_6n57), .CO(vscale_core_DW01_sub_6n56), .S(pipeline_md_N311) );
  FA_X1 vscale_core_DW01_sub_6_U5 ( .A(vscale_core_DW01_sub_6n403), .B(pipeline_md_a[59]), .CI(vscale_core_DW01_sub_6n58), .CO(vscale_core_DW01_sub_6n57), .S(pipeline_md_N310) );
  FA_X1 vscale_core_DW01_sub_6_U6 ( .A(vscale_core_DW01_sub_6n404), .B(pipeline_md_a[58]), .CI(vscale_core_DW01_sub_6n59), .CO(vscale_core_DW01_sub_6n58), .S(pipeline_md_N309) );
  FA_X1 vscale_core_DW01_sub_6_U7 ( .A(vscale_core_DW01_sub_6n405), .B(pipeline_md_a[57]), .CI(vscale_core_DW01_sub_6n60), .CO(vscale_core_DW01_sub_6n59), .S(pipeline_md_N308) );
  FA_X1 vscale_core_DW01_sub_6_U8 ( .A(vscale_core_DW01_sub_6n406), .B(pipeline_md_a[56]), .CI(vscale_core_DW01_sub_6n61), .CO(vscale_core_DW01_sub_6n60), .S(pipeline_md_N307) );
  FA_X1 vscale_core_DW01_sub_6_U9 ( .A(vscale_core_DW01_sub_6n407), .B(pipeline_md_a[55]), .CI(vscale_core_DW01_sub_6n62), .CO(vscale_core_DW01_sub_6n61), .S(pipeline_md_N306) );
  FA_X1 vscale_core_DW01_sub_6_U10 ( .A(vscale_core_DW01_sub_6n408), .B(pipeline_md_a[54]), .CI(vscale_core_DW01_sub_6n63), .CO(vscale_core_DW01_sub_6n62), .S(pipeline_md_N305) );
  XOR2_X2 vscale_core_DW01_sub_6_U11 ( .A(vscale_core_DW01_sub_6n1), .B(vscale_core_DW01_sub_6n66), .Z(pipeline_md_N304) );
  NAND2_X2 vscale_core_DW01_sub_6_U13 ( .A1(vscale_core_DW01_sub_6n347), .A2(vscale_core_DW01_sub_6n65), .ZN(vscale_core_DW01_sub_6n1) );
  NAND2_X2 vscale_core_DW01_sub_6_U16 ( .A1(vscale_core_DW01_sub_6n409), .A2(pipeline_md_a[53]), .ZN(vscale_core_DW01_sub_6n65) );
  XNOR2_X2 vscale_core_DW01_sub_6_U17 ( .A(vscale_core_DW01_sub_6n71), .B(vscale_core_DW01_sub_6n2), .ZN(pipeline_md_N303) );
  NAND2_X2 vscale_core_DW01_sub_6_U21 ( .A1(vscale_core_DW01_sub_6n665), .A2(vscale_core_DW01_sub_6n70), .ZN(vscale_core_DW01_sub_6n2) );
  NAND2_X2 vscale_core_DW01_sub_6_U24 ( .A1(vscale_core_DW01_sub_6n410), .A2(pipeline_md_a[52]), .ZN(vscale_core_DW01_sub_6n70) );
  XOR2_X2 vscale_core_DW01_sub_6_U25 ( .A(vscale_core_DW01_sub_6n3), .B(vscale_core_DW01_sub_6n74), .Z(pipeline_md_N302) );
  NAND2_X2 vscale_core_DW01_sub_6_U27 ( .A1(vscale_core_DW01_sub_6n349), .A2(vscale_core_DW01_sub_6n73), .ZN(vscale_core_DW01_sub_6n3) );
  NAND2_X2 vscale_core_DW01_sub_6_U30 ( .A1(vscale_core_DW01_sub_6n411), .A2(pipeline_md_a[51]), .ZN(vscale_core_DW01_sub_6n73) );
  XNOR2_X2 vscale_core_DW01_sub_6_U31 ( .A(vscale_core_DW01_sub_6n79), .B(vscale_core_DW01_sub_6n4), .ZN(pipeline_md_N301) );
  NAND2_X2 vscale_core_DW01_sub_6_U35 ( .A1(vscale_core_DW01_sub_6n664), .A2(vscale_core_DW01_sub_6n78), .ZN(vscale_core_DW01_sub_6n4) );
  NAND2_X2 vscale_core_DW01_sub_6_U38 ( .A1(vscale_core_DW01_sub_6n412), .A2(pipeline_md_a[50]), .ZN(vscale_core_DW01_sub_6n78) );
  XOR2_X2 vscale_core_DW01_sub_6_U39 ( .A(vscale_core_DW01_sub_6n5), .B(vscale_core_DW01_sub_6n82), .Z(pipeline_md_N300) );
  NAND2_X2 vscale_core_DW01_sub_6_U41 ( .A1(vscale_core_DW01_sub_6n351), .A2(vscale_core_DW01_sub_6n81), .ZN(vscale_core_DW01_sub_6n5) );
  NAND2_X2 vscale_core_DW01_sub_6_U44 ( .A1(vscale_core_DW01_sub_6n413), .A2(pipeline_md_a[49]), .ZN(vscale_core_DW01_sub_6n81) );
  XNOR2_X2 vscale_core_DW01_sub_6_U45 ( .A(vscale_core_DW01_sub_6n87), .B(vscale_core_DW01_sub_6n6), .ZN(pipeline_md_N299) );
  NAND2_X2 vscale_core_DW01_sub_6_U49 ( .A1(vscale_core_DW01_sub_6n662), .A2(vscale_core_DW01_sub_6n86), .ZN(vscale_core_DW01_sub_6n6) );
  NAND2_X2 vscale_core_DW01_sub_6_U52 ( .A1(vscale_core_DW01_sub_6n414), .A2(pipeline_md_a[48]), .ZN(vscale_core_DW01_sub_6n86) );
  XOR2_X2 vscale_core_DW01_sub_6_U53 ( .A(vscale_core_DW01_sub_6n7), .B(vscale_core_DW01_sub_6n90), .Z(pipeline_md_N298) );
  NAND2_X2 vscale_core_DW01_sub_6_U55 ( .A1(vscale_core_DW01_sub_6n353), .A2(vscale_core_DW01_sub_6n89), .ZN(vscale_core_DW01_sub_6n7) );
  NAND2_X2 vscale_core_DW01_sub_6_U58 ( .A1(vscale_core_DW01_sub_6n415), .A2(pipeline_md_a[47]), .ZN(vscale_core_DW01_sub_6n89) );
  XNOR2_X2 vscale_core_DW01_sub_6_U59 ( .A(vscale_core_DW01_sub_6n95), .B(vscale_core_DW01_sub_6n8), .ZN(pipeline_md_N297) );
  NAND2_X2 vscale_core_DW01_sub_6_U63 ( .A1(vscale_core_DW01_sub_6n661), .A2(vscale_core_DW01_sub_6n94), .ZN(vscale_core_DW01_sub_6n8) );
  NAND2_X2 vscale_core_DW01_sub_6_U66 ( .A1(vscale_core_DW01_sub_6n416), .A2(pipeline_md_a[46]), .ZN(vscale_core_DW01_sub_6n94) );
  XOR2_X2 vscale_core_DW01_sub_6_U67 ( .A(vscale_core_DW01_sub_6n9), .B(vscale_core_DW01_sub_6n98), .Z(pipeline_md_N296) );
  NAND2_X2 vscale_core_DW01_sub_6_U69 ( .A1(vscale_core_DW01_sub_6n355), .A2(vscale_core_DW01_sub_6n97), .ZN(vscale_core_DW01_sub_6n9) );
  NAND2_X2 vscale_core_DW01_sub_6_U72 ( .A1(vscale_core_DW01_sub_6n417), .A2(pipeline_md_a[45]), .ZN(vscale_core_DW01_sub_6n97) );
  XNOR2_X2 vscale_core_DW01_sub_6_U73 ( .A(vscale_core_DW01_sub_6n103), .B(vscale_core_DW01_sub_6n10), .ZN(pipeline_md_N295) );
  NAND2_X2 vscale_core_DW01_sub_6_U77 ( .A1(vscale_core_DW01_sub_6n663), .A2(vscale_core_DW01_sub_6n102), .ZN(vscale_core_DW01_sub_6n10) );
  NAND2_X2 vscale_core_DW01_sub_6_U80 ( .A1(vscale_core_DW01_sub_6n418), .A2(pipeline_md_a[44]), .ZN(vscale_core_DW01_sub_6n102) );
  XOR2_X2 vscale_core_DW01_sub_6_U81 ( .A(vscale_core_DW01_sub_6n11), .B(vscale_core_DW01_sub_6n106), .Z(pipeline_md_N294) );
  NAND2_X2 vscale_core_DW01_sub_6_U83 ( .A1(vscale_core_DW01_sub_6n357), .A2(vscale_core_DW01_sub_6n105), .ZN(vscale_core_DW01_sub_6n11) );
  NAND2_X2 vscale_core_DW01_sub_6_U86 ( .A1(vscale_core_DW01_sub_6n419), .A2(pipeline_md_a[43]), .ZN(vscale_core_DW01_sub_6n105) );
  XNOR2_X2 vscale_core_DW01_sub_6_U87 ( .A(vscale_core_DW01_sub_6n111), .B(vscale_core_DW01_sub_6n12), .ZN(pipeline_md_N293) );
  NAND2_X2 vscale_core_DW01_sub_6_U91 ( .A1(vscale_core_DW01_sub_6n358), .A2(vscale_core_DW01_sub_6n110), .ZN(vscale_core_DW01_sub_6n12) );
  NAND2_X2 vscale_core_DW01_sub_6_U94 ( .A1(vscale_core_DW01_sub_6n420), .A2(pipeline_md_a[42]), .ZN(vscale_core_DW01_sub_6n110) );
  XOR2_X2 vscale_core_DW01_sub_6_U95 ( .A(vscale_core_DW01_sub_6n13), .B(vscale_core_DW01_sub_6n118), .Z(pipeline_md_N292) );
  NAND2_X2 vscale_core_DW01_sub_6_U97 ( .A1(vscale_core_DW01_sub_6n126), .A2(vscale_core_DW01_sub_6n114), .ZN(vscale_core_DW01_sub_6n112) );
  NAND2_X2 vscale_core_DW01_sub_6_U101 ( .A1(vscale_core_DW01_sub_6n359), .A2(vscale_core_DW01_sub_6n117), .ZN(vscale_core_DW01_sub_6n13) );
  NAND2_X2 vscale_core_DW01_sub_6_U104 ( .A1(vscale_core_DW01_sub_6n421), .A2(pipeline_md_a[41]), .ZN(vscale_core_DW01_sub_6n117) );
  XNOR2_X2 vscale_core_DW01_sub_6_U105 ( .A(vscale_core_DW01_sub_6n123), .B(vscale_core_DW01_sub_6n14), .ZN(pipeline_md_N291) );
  NAND2_X2 vscale_core_DW01_sub_6_U109 ( .A1(vscale_core_DW01_sub_6n360), .A2(vscale_core_DW01_sub_6n122), .ZN(vscale_core_DW01_sub_6n14) );
  NAND2_X2 vscale_core_DW01_sub_6_U112 ( .A1(vscale_core_DW01_sub_6n422), .A2(pipeline_md_a[40]), .ZN(vscale_core_DW01_sub_6n122) );
  XOR2_X2 vscale_core_DW01_sub_6_U113 ( .A(vscale_core_DW01_sub_6n15), .B(vscale_core_DW01_sub_6n134), .Z(pipeline_md_N290) );
  NAND2_X2 vscale_core_DW01_sub_6_U119 ( .A1(vscale_core_DW01_sub_6n142), .A2(vscale_core_DW01_sub_6n130), .ZN(vscale_core_DW01_sub_6n128) );
  NAND2_X2 vscale_core_DW01_sub_6_U123 ( .A1(vscale_core_DW01_sub_6n361), .A2(vscale_core_DW01_sub_6n133), .ZN(vscale_core_DW01_sub_6n15) );
  NAND2_X2 vscale_core_DW01_sub_6_U126 ( .A1(vscale_core_DW01_sub_6n423), .A2(pipeline_md_a[39]), .ZN(vscale_core_DW01_sub_6n133) );
  XNOR2_X2 vscale_core_DW01_sub_6_U127 ( .A(vscale_core_DW01_sub_6n139), .B(vscale_core_DW01_sub_6n16), .ZN(pipeline_md_N289) );
  NAND2_X2 vscale_core_DW01_sub_6_U131 ( .A1(vscale_core_DW01_sub_6n362), .A2(vscale_core_DW01_sub_6n138), .ZN(vscale_core_DW01_sub_6n16) );
  NAND2_X2 vscale_core_DW01_sub_6_U134 ( .A1(vscale_core_DW01_sub_6n424), .A2(pipeline_md_a[38]), .ZN(vscale_core_DW01_sub_6n138) );
  XOR2_X2 vscale_core_DW01_sub_6_U135 ( .A(vscale_core_DW01_sub_6n17), .B(vscale_core_DW01_sub_6n146), .Z(pipeline_md_N288) );
  NAND2_X2 vscale_core_DW01_sub_6_U141 ( .A1(vscale_core_DW01_sub_6n363), .A2(vscale_core_DW01_sub_6n145), .ZN(vscale_core_DW01_sub_6n17) );
  NAND2_X2 vscale_core_DW01_sub_6_U144 ( .A1(vscale_core_DW01_sub_6n425), .A2(pipeline_md_a[37]), .ZN(vscale_core_DW01_sub_6n145) );
  XOR2_X2 vscale_core_DW01_sub_6_U145 ( .A(vscale_core_DW01_sub_6n18), .B(vscale_core_DW01_sub_6n151), .Z(pipeline_md_N287) );
  NAND2_X2 vscale_core_DW01_sub_6_U149 ( .A1(vscale_core_DW01_sub_6n364), .A2(vscale_core_DW01_sub_6n150), .ZN(vscale_core_DW01_sub_6n18) );
  NAND2_X2 vscale_core_DW01_sub_6_U152 ( .A1(vscale_core_DW01_sub_6n426), .A2(pipeline_md_a[36]), .ZN(vscale_core_DW01_sub_6n150) );
  XOR2_X2 vscale_core_DW01_sub_6_U153 ( .A(vscale_core_DW01_sub_6n19), .B(vscale_core_DW01_sub_6n159), .Z(pipeline_md_N286) );
  NAND2_X2 vscale_core_DW01_sub_6_U156 ( .A1(vscale_core_DW01_sub_6n167), .A2(vscale_core_DW01_sub_6n155), .ZN(vscale_core_DW01_sub_6n153) );
  NAND2_X2 vscale_core_DW01_sub_6_U160 ( .A1(vscale_core_DW01_sub_6n365), .A2(vscale_core_DW01_sub_6n158), .ZN(vscale_core_DW01_sub_6n19) );
  NAND2_X2 vscale_core_DW01_sub_6_U163 ( .A1(vscale_core_DW01_sub_6n427), .A2(pipeline_md_a[35]), .ZN(vscale_core_DW01_sub_6n158) );
  XNOR2_X2 vscale_core_DW01_sub_6_U164 ( .A(vscale_core_DW01_sub_6n164), .B(vscale_core_DW01_sub_6n20), .ZN(pipeline_md_N285) );
  NAND2_X2 vscale_core_DW01_sub_6_U168 ( .A1(vscale_core_DW01_sub_6n366), .A2(vscale_core_DW01_sub_6n163), .ZN(vscale_core_DW01_sub_6n20) );
  NAND2_X2 vscale_core_DW01_sub_6_U171 ( .A1(vscale_core_DW01_sub_6n428), .A2(pipeline_md_a[34]), .ZN(vscale_core_DW01_sub_6n163) );
  XNOR2_X2 vscale_core_DW01_sub_6_U172 ( .A(vscale_core_DW01_sub_6n171), .B(vscale_core_DW01_sub_6n21), .ZN(pipeline_md_N284) );
  NAND2_X2 vscale_core_DW01_sub_6_U178 ( .A1(vscale_core_DW01_sub_6n367), .A2(vscale_core_DW01_sub_6n170), .ZN(vscale_core_DW01_sub_6n21) );
  NAND2_X2 vscale_core_DW01_sub_6_U181 ( .A1(vscale_core_DW01_sub_6n429), .A2(pipeline_md_a[33]), .ZN(vscale_core_DW01_sub_6n170) );
  XOR2_X2 vscale_core_DW01_sub_6_U182 ( .A(vscale_core_DW01_sub_6n22), .B(vscale_core_DW01_sub_6n174), .Z(pipeline_md_N283) );
  NAND2_X2 vscale_core_DW01_sub_6_U184 ( .A1(vscale_core_DW01_sub_6n368), .A2(vscale_core_DW01_sub_6n173), .ZN(vscale_core_DW01_sub_6n22) );
  NAND2_X2 vscale_core_DW01_sub_6_U187 ( .A1(vscale_core_DW01_sub_6n430), .A2(pipeline_md_a[32]), .ZN(vscale_core_DW01_sub_6n173) );
  XNOR2_X2 vscale_core_DW01_sub_6_U188 ( .A(vscale_core_DW01_sub_6n186), .B(vscale_core_DW01_sub_6n23), .ZN(pipeline_md_N282) );
  NAND2_X2 vscale_core_DW01_sub_6_U191 ( .A1(vscale_core_DW01_sub_6n220), .A2(vscale_core_DW01_sub_6n178), .ZN(vscale_core_DW01_sub_6n176) );
  NAND2_X2 vscale_core_DW01_sub_6_U195 ( .A1(vscale_core_DW01_sub_6n190), .A2(vscale_core_DW01_sub_6n182), .ZN(vscale_core_DW01_sub_6n180) );
  NAND2_X2 vscale_core_DW01_sub_6_U199 ( .A1(vscale_core_DW01_sub_6n369), .A2(vscale_core_DW01_sub_6n185), .ZN(vscale_core_DW01_sub_6n23) );
  NAND2_X2 vscale_core_DW01_sub_6_U202 ( .A1(vscale_core_DW01_sub_6n431), .A2(pipeline_md_a[31]), .ZN(vscale_core_DW01_sub_6n185) );
  XOR2_X2 vscale_core_DW01_sub_6_U203 ( .A(vscale_core_DW01_sub_6n24), .B(vscale_core_DW01_sub_6n189), .Z(pipeline_md_N281) );
  NAND2_X2 vscale_core_DW01_sub_6_U205 ( .A1(vscale_core_DW01_sub_6n370), .A2(vscale_core_DW01_sub_6n188), .ZN(vscale_core_DW01_sub_6n24) );
  NAND2_X2 vscale_core_DW01_sub_6_U208 ( .A1(vscale_core_DW01_sub_6n432), .A2(pipeline_md_a[30]), .ZN(vscale_core_DW01_sub_6n188) );
  XNOR2_X2 vscale_core_DW01_sub_6_U209 ( .A(vscale_core_DW01_sub_6n194), .B(vscale_core_DW01_sub_6n25), .ZN(pipeline_md_N280) );
  NAND2_X2 vscale_core_DW01_sub_6_U213 ( .A1(vscale_core_DW01_sub_6n371), .A2(vscale_core_DW01_sub_6n193), .ZN(vscale_core_DW01_sub_6n25) );
  NAND2_X2 vscale_core_DW01_sub_6_U216 ( .A1(vscale_core_DW01_sub_6n433), .A2(pipeline_md_a[29]), .ZN(vscale_core_DW01_sub_6n193) );
  XNOR2_X2 vscale_core_DW01_sub_6_U217 ( .A(vscale_core_DW01_sub_6n197), .B(vscale_core_DW01_sub_6n26), .ZN(pipeline_md_N279) );
  NAND2_X2 vscale_core_DW01_sub_6_U219 ( .A1(vscale_core_DW01_sub_6n372), .A2(vscale_core_DW01_sub_6n196), .ZN(vscale_core_DW01_sub_6n26) );
  NAND2_X2 vscale_core_DW01_sub_6_U222 ( .A1(vscale_core_DW01_sub_6n434), .A2(pipeline_md_a[28]), .ZN(vscale_core_DW01_sub_6n196) );
  XNOR2_X2 vscale_core_DW01_sub_6_U223 ( .A(vscale_core_DW01_sub_6n207), .B(vscale_core_DW01_sub_6n27), .ZN(pipeline_md_N278) );
  NAND2_X2 vscale_core_DW01_sub_6_U228 ( .A1(vscale_core_DW01_sub_6n211), .A2(vscale_core_DW01_sub_6n203), .ZN(vscale_core_DW01_sub_6n201) );
  NAND2_X2 vscale_core_DW01_sub_6_U232 ( .A1(vscale_core_DW01_sub_6n373), .A2(vscale_core_DW01_sub_6n206), .ZN(vscale_core_DW01_sub_6n27) );
  NAND2_X2 vscale_core_DW01_sub_6_U235 ( .A1(vscale_core_DW01_sub_6n435), .A2(pipeline_md_a[27]), .ZN(vscale_core_DW01_sub_6n206) );
  XOR2_X2 vscale_core_DW01_sub_6_U236 ( .A(vscale_core_DW01_sub_6n28), .B(vscale_core_DW01_sub_6n210), .Z(pipeline_md_N277) );
  NAND2_X2 vscale_core_DW01_sub_6_U238 ( .A1(vscale_core_DW01_sub_6n374), .A2(vscale_core_DW01_sub_6n209), .ZN(vscale_core_DW01_sub_6n28) );
  NAND2_X2 vscale_core_DW01_sub_6_U241 ( .A1(vscale_core_DW01_sub_6n436), .A2(pipeline_md_a[26]), .ZN(vscale_core_DW01_sub_6n209) );
  XNOR2_X2 vscale_core_DW01_sub_6_U242 ( .A(vscale_core_DW01_sub_6n215), .B(vscale_core_DW01_sub_6n29), .ZN(pipeline_md_N276) );
  NAND2_X2 vscale_core_DW01_sub_6_U246 ( .A1(vscale_core_DW01_sub_6n375), .A2(vscale_core_DW01_sub_6n214), .ZN(vscale_core_DW01_sub_6n29) );
  NAND2_X2 vscale_core_DW01_sub_6_U249 ( .A1(vscale_core_DW01_sub_6n437), .A2(pipeline_md_a[25]), .ZN(vscale_core_DW01_sub_6n214) );
  XNOR2_X2 vscale_core_DW01_sub_6_U250 ( .A(vscale_core_DW01_sub_6n218), .B(vscale_core_DW01_sub_6n30), .ZN(pipeline_md_N275) );
  NAND2_X2 vscale_core_DW01_sub_6_U252 ( .A1(vscale_core_DW01_sub_6n376), .A2(vscale_core_DW01_sub_6n217), .ZN(vscale_core_DW01_sub_6n30) );
  NAND2_X2 vscale_core_DW01_sub_6_U255 ( .A1(vscale_core_DW01_sub_6n438), .A2(pipeline_md_a[24]), .ZN(vscale_core_DW01_sub_6n217) );
  XNOR2_X2 vscale_core_DW01_sub_6_U256 ( .A(vscale_core_DW01_sub_6n228), .B(vscale_core_DW01_sub_6n31), .ZN(pipeline_md_N274) );
  NAND2_X2 vscale_core_DW01_sub_6_U261 ( .A1(vscale_core_DW01_sub_6n232), .A2(vscale_core_DW01_sub_6n224), .ZN(vscale_core_DW01_sub_6n222) );
  NAND2_X2 vscale_core_DW01_sub_6_U265 ( .A1(vscale_core_DW01_sub_6n377), .A2(vscale_core_DW01_sub_6n227), .ZN(vscale_core_DW01_sub_6n31) );
  NAND2_X2 vscale_core_DW01_sub_6_U268 ( .A1(vscale_core_DW01_sub_6n439), .A2(pipeline_md_a[23]), .ZN(vscale_core_DW01_sub_6n227) );
  XOR2_X2 vscale_core_DW01_sub_6_U269 ( .A(vscale_core_DW01_sub_6n32), .B(vscale_core_DW01_sub_6n231), .Z(pipeline_md_N273) );
  NAND2_X2 vscale_core_DW01_sub_6_U271 ( .A1(vscale_core_DW01_sub_6n378), .A2(vscale_core_DW01_sub_6n230), .ZN(vscale_core_DW01_sub_6n32) );
  NAND2_X2 vscale_core_DW01_sub_6_U274 ( .A1(vscale_core_DW01_sub_6n440), .A2(pipeline_md_a[22]), .ZN(vscale_core_DW01_sub_6n230) );
  XNOR2_X2 vscale_core_DW01_sub_6_U275 ( .A(vscale_core_DW01_sub_6n236), .B(vscale_core_DW01_sub_6n33), .ZN(pipeline_md_N272) );
  NAND2_X2 vscale_core_DW01_sub_6_U279 ( .A1(vscale_core_DW01_sub_6n379), .A2(vscale_core_DW01_sub_6n235), .ZN(vscale_core_DW01_sub_6n33) );
  NAND2_X2 vscale_core_DW01_sub_6_U282 ( .A1(vscale_core_DW01_sub_6n441), .A2(pipeline_md_a[21]), .ZN(vscale_core_DW01_sub_6n235) );
  XNOR2_X2 vscale_core_DW01_sub_6_U283 ( .A(vscale_core_DW01_sub_6n239), .B(vscale_core_DW01_sub_6n34), .ZN(pipeline_md_N271) );
  NAND2_X2 vscale_core_DW01_sub_6_U285 ( .A1(vscale_core_DW01_sub_6n380), .A2(vscale_core_DW01_sub_6n238), .ZN(vscale_core_DW01_sub_6n34) );
  NAND2_X2 vscale_core_DW01_sub_6_U288 ( .A1(vscale_core_DW01_sub_6n442), .A2(pipeline_md_a[20]), .ZN(vscale_core_DW01_sub_6n238) );
  XNOR2_X2 vscale_core_DW01_sub_6_U289 ( .A(vscale_core_DW01_sub_6n249), .B(vscale_core_DW01_sub_6n35), .ZN(pipeline_md_N270) );
  NAND2_X2 vscale_core_DW01_sub_6_U294 ( .A1(vscale_core_DW01_sub_6n253), .A2(vscale_core_DW01_sub_6n245), .ZN(vscale_core_DW01_sub_6n243) );
  NAND2_X2 vscale_core_DW01_sub_6_U298 ( .A1(vscale_core_DW01_sub_6n381), .A2(vscale_core_DW01_sub_6n248), .ZN(vscale_core_DW01_sub_6n35) );
  NAND2_X2 vscale_core_DW01_sub_6_U301 ( .A1(vscale_core_DW01_sub_6n443), .A2(pipeline_md_a[19]), .ZN(vscale_core_DW01_sub_6n248) );
  XOR2_X2 vscale_core_DW01_sub_6_U302 ( .A(vscale_core_DW01_sub_6n36), .B(vscale_core_DW01_sub_6n252), .Z(pipeline_md_N269) );
  NAND2_X2 vscale_core_DW01_sub_6_U304 ( .A1(vscale_core_DW01_sub_6n382), .A2(vscale_core_DW01_sub_6n251), .ZN(vscale_core_DW01_sub_6n36) );
  NAND2_X2 vscale_core_DW01_sub_6_U307 ( .A1(vscale_core_DW01_sub_6n444), .A2(pipeline_md_a[18]), .ZN(vscale_core_DW01_sub_6n251) );
  XOR2_X2 vscale_core_DW01_sub_6_U308 ( .A(vscale_core_DW01_sub_6n37), .B(vscale_core_DW01_sub_6n257), .Z(pipeline_md_N268) );
  NAND2_X2 vscale_core_DW01_sub_6_U312 ( .A1(vscale_core_DW01_sub_6n383), .A2(vscale_core_DW01_sub_6n256), .ZN(vscale_core_DW01_sub_6n37) );
  NAND2_X2 vscale_core_DW01_sub_6_U315 ( .A1(vscale_core_DW01_sub_6n445), .A2(pipeline_md_a[17]), .ZN(vscale_core_DW01_sub_6n256) );
  XNOR2_X2 vscale_core_DW01_sub_6_U316 ( .A(vscale_core_DW01_sub_6n262), .B(vscale_core_DW01_sub_6n38), .ZN(pipeline_md_N267) );
  NAND2_X2 vscale_core_DW01_sub_6_U320 ( .A1(vscale_core_DW01_sub_6n384), .A2(vscale_core_DW01_sub_6n261), .ZN(vscale_core_DW01_sub_6n38) );
  NAND2_X2 vscale_core_DW01_sub_6_U323 ( .A1(vscale_core_DW01_sub_6n446), .A2(pipeline_md_a[16]), .ZN(vscale_core_DW01_sub_6n261) );
  XOR2_X2 vscale_core_DW01_sub_6_U324 ( .A(vscale_core_DW01_sub_6n39), .B(vscale_core_DW01_sub_6n272), .Z(pipeline_md_N266) );
  NAND2_X2 vscale_core_DW01_sub_6_U329 ( .A1(vscale_core_DW01_sub_6n280), .A2(vscale_core_DW01_sub_6n268), .ZN(vscale_core_DW01_sub_6n266) );
  NAND2_X2 vscale_core_DW01_sub_6_U333 ( .A1(vscale_core_DW01_sub_6n385), .A2(vscale_core_DW01_sub_6n271), .ZN(vscale_core_DW01_sub_6n39) );
  NAND2_X2 vscale_core_DW01_sub_6_U336 ( .A1(vscale_core_DW01_sub_6n447), .A2(pipeline_md_a[15]), .ZN(vscale_core_DW01_sub_6n271) );
  XNOR2_X2 vscale_core_DW01_sub_6_U337 ( .A(vscale_core_DW01_sub_6n277), .B(vscale_core_DW01_sub_6n40), .ZN(pipeline_md_N265) );
  NAND2_X2 vscale_core_DW01_sub_6_U341 ( .A1(vscale_core_DW01_sub_6n386), .A2(vscale_core_DW01_sub_6n276), .ZN(vscale_core_DW01_sub_6n40) );
  NAND2_X2 vscale_core_DW01_sub_6_U344 ( .A1(vscale_core_DW01_sub_6n448), .A2(pipeline_md_a[14]), .ZN(vscale_core_DW01_sub_6n276) );
  XOR2_X2 vscale_core_DW01_sub_6_U345 ( .A(vscale_core_DW01_sub_6n41), .B(vscale_core_DW01_sub_6n284), .Z(pipeline_md_N264) );
  NAND2_X2 vscale_core_DW01_sub_6_U351 ( .A1(vscale_core_DW01_sub_6n387), .A2(vscale_core_DW01_sub_6n283), .ZN(vscale_core_DW01_sub_6n41) );
  NAND2_X2 vscale_core_DW01_sub_6_U354 ( .A1(vscale_core_DW01_sub_6n449), .A2(pipeline_md_a[13]), .ZN(vscale_core_DW01_sub_6n283) );
  XOR2_X2 vscale_core_DW01_sub_6_U355 ( .A(vscale_core_DW01_sub_6n42), .B(vscale_core_DW01_sub_6n289), .Z(pipeline_md_N263) );
  NAND2_X2 vscale_core_DW01_sub_6_U359 ( .A1(vscale_core_DW01_sub_6n388), .A2(vscale_core_DW01_sub_6n288), .ZN(vscale_core_DW01_sub_6n42) );
  NAND2_X2 vscale_core_DW01_sub_6_U362 ( .A1(vscale_core_DW01_sub_6n450), .A2(pipeline_md_a[12]), .ZN(vscale_core_DW01_sub_6n288) );
  XOR2_X2 vscale_core_DW01_sub_6_U363 ( .A(vscale_core_DW01_sub_6n43), .B(vscale_core_DW01_sub_6n297), .Z(pipeline_md_N262) );
  NAND2_X2 vscale_core_DW01_sub_6_U366 ( .A1(vscale_core_DW01_sub_6n305), .A2(vscale_core_DW01_sub_6n293), .ZN(vscale_core_DW01_sub_6n291) );
  NAND2_X2 vscale_core_DW01_sub_6_U370 ( .A1(vscale_core_DW01_sub_6n389), .A2(vscale_core_DW01_sub_6n296), .ZN(vscale_core_DW01_sub_6n43) );
  NAND2_X2 vscale_core_DW01_sub_6_U373 ( .A1(vscale_core_DW01_sub_6n451), .A2(pipeline_md_a[11]), .ZN(vscale_core_DW01_sub_6n296) );
  XNOR2_X2 vscale_core_DW01_sub_6_U374 ( .A(vscale_core_DW01_sub_6n302), .B(vscale_core_DW01_sub_6n44), .ZN(pipeline_md_N261) );
  NAND2_X2 vscale_core_DW01_sub_6_U378 ( .A1(vscale_core_DW01_sub_6n390), .A2(vscale_core_DW01_sub_6n301), .ZN(vscale_core_DW01_sub_6n44) );
  NAND2_X2 vscale_core_DW01_sub_6_U381 ( .A1(vscale_core_DW01_sub_6n452), .A2(pipeline_md_a[10]), .ZN(vscale_core_DW01_sub_6n301) );
  XNOR2_X2 vscale_core_DW01_sub_6_U382 ( .A(vscale_core_DW01_sub_6n309), .B(vscale_core_DW01_sub_6n45), .ZN(pipeline_md_N260) );
  NAND2_X2 vscale_core_DW01_sub_6_U388 ( .A1(vscale_core_DW01_sub_6n391), .A2(vscale_core_DW01_sub_6n308), .ZN(vscale_core_DW01_sub_6n45) );
  NAND2_X2 vscale_core_DW01_sub_6_U391 ( .A1(vscale_core_DW01_sub_6n453), .A2(pipeline_md_a[9]), .ZN(vscale_core_DW01_sub_6n308) );
  XOR2_X2 vscale_core_DW01_sub_6_U392 ( .A(vscale_core_DW01_sub_6n46), .B(vscale_core_DW01_sub_6n312), .Z(pipeline_md_N259) );
  NAND2_X2 vscale_core_DW01_sub_6_U394 ( .A1(vscale_core_DW01_sub_6n392), .A2(vscale_core_DW01_sub_6n311), .ZN(vscale_core_DW01_sub_6n46) );
  NAND2_X2 vscale_core_DW01_sub_6_U397 ( .A1(vscale_core_DW01_sub_6n454), .A2(pipeline_md_a[8]), .ZN(vscale_core_DW01_sub_6n311) );
  XNOR2_X2 vscale_core_DW01_sub_6_U398 ( .A(vscale_core_DW01_sub_6n320), .B(vscale_core_DW01_sub_6n47), .ZN(pipeline_md_N258) );
  NAND2_X2 vscale_core_DW01_sub_6_U401 ( .A1(vscale_core_DW01_sub_6n324), .A2(vscale_core_DW01_sub_6n316), .ZN(vscale_core_DW01_sub_6n314) );
  NAND2_X2 vscale_core_DW01_sub_6_U405 ( .A1(vscale_core_DW01_sub_6n393), .A2(vscale_core_DW01_sub_6n319), .ZN(vscale_core_DW01_sub_6n47) );
  NAND2_X2 vscale_core_DW01_sub_6_U408 ( .A1(vscale_core_DW01_sub_6n455), .A2(pipeline_md_a[7]), .ZN(vscale_core_DW01_sub_6n319) );
  XOR2_X2 vscale_core_DW01_sub_6_U409 ( .A(vscale_core_DW01_sub_6n48), .B(vscale_core_DW01_sub_6n323), .Z(pipeline_md_N257) );
  NAND2_X2 vscale_core_DW01_sub_6_U411 ( .A1(vscale_core_DW01_sub_6n394), .A2(vscale_core_DW01_sub_6n322), .ZN(vscale_core_DW01_sub_6n48) );
  NAND2_X2 vscale_core_DW01_sub_6_U414 ( .A1(vscale_core_DW01_sub_6n456), .A2(pipeline_md_a[6]), .ZN(vscale_core_DW01_sub_6n322) );
  XOR2_X2 vscale_core_DW01_sub_6_U415 ( .A(vscale_core_DW01_sub_6n49), .B(vscale_core_DW01_sub_6n328), .Z(pipeline_md_N256) );
  NAND2_X2 vscale_core_DW01_sub_6_U419 ( .A1(vscale_core_DW01_sub_6n395), .A2(vscale_core_DW01_sub_6n327), .ZN(vscale_core_DW01_sub_6n49) );
  NAND2_X2 vscale_core_DW01_sub_6_U422 ( .A1(vscale_core_DW01_sub_6n457), .A2(pipeline_md_a[5]), .ZN(vscale_core_DW01_sub_6n327) );
  XNOR2_X2 vscale_core_DW01_sub_6_U423 ( .A(vscale_core_DW01_sub_6n333), .B(vscale_core_DW01_sub_6n50), .ZN(pipeline_md_N255) );
  NAND2_X2 vscale_core_DW01_sub_6_U427 ( .A1(vscale_core_DW01_sub_6n396), .A2(vscale_core_DW01_sub_6n332), .ZN(vscale_core_DW01_sub_6n50) );
  NAND2_X2 vscale_core_DW01_sub_6_U430 ( .A1(vscale_core_DW01_sub_6n458), .A2(pipeline_md_a[4]), .ZN(vscale_core_DW01_sub_6n332) );
  XNOR2_X2 vscale_core_DW01_sub_6_U431 ( .A(vscale_core_DW01_sub_6n339), .B(vscale_core_DW01_sub_6n51), .ZN(pipeline_md_N254) );
  NAND2_X2 vscale_core_DW01_sub_6_U436 ( .A1(vscale_core_DW01_sub_6n397), .A2(vscale_core_DW01_sub_6n338), .ZN(vscale_core_DW01_sub_6n51) );
  NAND2_X2 vscale_core_DW01_sub_6_U439 ( .A1(vscale_core_DW01_sub_6n459), .A2(pipeline_md_a[3]), .ZN(vscale_core_DW01_sub_6n338) );
  XOR2_X2 vscale_core_DW01_sub_6_U440 ( .A(vscale_core_DW01_sub_6n52), .B(vscale_core_DW01_sub_6n342), .Z(pipeline_md_N253) );
  NAND2_X2 vscale_core_DW01_sub_6_U442 ( .A1(vscale_core_DW01_sub_6n398), .A2(vscale_core_DW01_sub_6n341), .ZN(vscale_core_DW01_sub_6n52) );
  NAND2_X2 vscale_core_DW01_sub_6_U445 ( .A1(vscale_core_DW01_sub_6n460), .A2(pipeline_md_a[2]), .ZN(vscale_core_DW01_sub_6n341) );
  XOR2_X2 vscale_core_DW01_sub_6_U446 ( .A(vscale_core_DW01_sub_6n346), .B(vscale_core_DW01_sub_6n53), .Z(pipeline_md_N252) );
  NAND2_X2 vscale_core_DW01_sub_6_U449 ( .A1(vscale_core_DW01_sub_6n399), .A2(vscale_core_DW01_sub_6n345), .ZN(vscale_core_DW01_sub_6n53) );
  NAND2_X2 vscale_core_DW01_sub_6_U452 ( .A1(vscale_core_DW01_sub_6n461), .A2(pipeline_md_a[1]), .ZN(vscale_core_DW01_sub_6n345) );
  XNOR2_X2 vscale_core_DW01_sub_6_U453 ( .A(vscale_core_DW01_sub_6n462), .B(pipeline_md_a[0]), .ZN(pipeline_md_N251) );
  NOR2_X2 vscale_core_DW01_sub_6_U521 ( .A1(vscale_core_DW01_sub_6n243), .A2(vscale_core_DW01_sub_6n222), .ZN(vscale_core_DW01_sub_6n220) );
  NOR2_X2 vscale_core_DW01_sub_6_U522 ( .A1(vscale_core_DW01_sub_6n153), .A2(vscale_core_DW01_sub_6n128), .ZN(vscale_core_DW01_sub_6n126) );
  AOI21_X2 vscale_core_DW01_sub_6_U523 ( .B1(vscale_core_DW01_sub_6n313), .B2(vscale_core_DW01_sub_6n264), .A(vscale_core_DW01_sub_6n265), .ZN(vscale_core_DW01_sub_6n263) );
  NOR2_X2 vscale_core_DW01_sub_6_U524 ( .A1(vscale_core_DW01_sub_6n291), .A2(vscale_core_DW01_sub_6n266), .ZN(vscale_core_DW01_sub_6n264) );
  OAI21_X2 vscale_core_DW01_sub_6_U525 ( .B1(vscale_core_DW01_sub_6n292), .B2(vscale_core_DW01_sub_6n266), .A(vscale_core_DW01_sub_6n267), .ZN(vscale_core_DW01_sub_6n265) );
  OAI21_X2 vscale_core_DW01_sub_6_U526 ( .B1(vscale_core_DW01_sub_6n263), .B2(vscale_core_DW01_sub_6n176), .A(vscale_core_DW01_sub_6n177), .ZN(vscale_core_DW01_sub_6n175) );
  AOI21_X2 vscale_core_DW01_sub_6_U527 ( .B1(vscale_core_DW01_sub_6n221), .B2(vscale_core_DW01_sub_6n178), .A(vscale_core_DW01_sub_6n179), .ZN(vscale_core_DW01_sub_6n177) );
  NOR2_X2 vscale_core_DW01_sub_6_U528 ( .A1(vscale_core_DW01_sub_6n201), .A2(vscale_core_DW01_sub_6n180), .ZN(vscale_core_DW01_sub_6n178) );
  AOI21_X2 vscale_core_DW01_sub_6_U529 ( .B1(vscale_core_DW01_sub_6n197), .B2(vscale_core_DW01_sub_6n190), .A(vscale_core_DW01_sub_6n191), .ZN(vscale_core_DW01_sub_6n189) );
  AOI21_X2 vscale_core_DW01_sub_6_U530 ( .B1(vscale_core_DW01_sub_6n218), .B2(vscale_core_DW01_sub_6n199), .A(vscale_core_DW01_sub_6n200), .ZN(vscale_core_DW01_sub_6n198) );
  AOI21_X2 vscale_core_DW01_sub_6_U531 ( .B1(vscale_core_DW01_sub_6n262), .B2(vscale_core_DW01_sub_6n220), .A(vscale_core_DW01_sub_6n221), .ZN(vscale_core_DW01_sub_6n219) );
  AOI21_X2 vscale_core_DW01_sub_6_U532 ( .B1(vscale_core_DW01_sub_6n218), .B2(vscale_core_DW01_sub_6n211), .A(vscale_core_DW01_sub_6n212), .ZN(vscale_core_DW01_sub_6n210) );
  AOI21_X2 vscale_core_DW01_sub_6_U533 ( .B1(vscale_core_DW01_sub_6n239), .B2(vscale_core_DW01_sub_6n232), .A(vscale_core_DW01_sub_6n233), .ZN(vscale_core_DW01_sub_6n231) );
  AOI21_X2 vscale_core_DW01_sub_6_U534 ( .B1(vscale_core_DW01_sub_6n262), .B2(vscale_core_DW01_sub_6n253), .A(vscale_core_DW01_sub_6n254), .ZN(vscale_core_DW01_sub_6n252) );
  AOI21_X2 vscale_core_DW01_sub_6_U535 ( .B1(vscale_core_DW01_sub_6n333), .B2(vscale_core_DW01_sub_6n324), .A(vscale_core_DW01_sub_6n325), .ZN(vscale_core_DW01_sub_6n323) );
  AOI21_X2 vscale_core_DW01_sub_6_U536 ( .B1(vscale_core_DW01_sub_6n262), .B2(vscale_core_DW01_sub_6n241), .A(vscale_core_DW01_sub_6n242), .ZN(vscale_core_DW01_sub_6n240) );
  OAI21_X2 vscale_core_DW01_sub_6_U537 ( .B1(vscale_core_DW01_sub_6n312), .B2(vscale_core_DW01_sub_6n291), .A(vscale_core_DW01_sub_6n292), .ZN(vscale_core_DW01_sub_6n290) );
  OAI21_X2 vscale_core_DW01_sub_6_U538 ( .B1(vscale_core_DW01_sub_6n174), .B2(vscale_core_DW01_sub_6n153), .A(vscale_core_DW01_sub_6n154), .ZN(vscale_core_DW01_sub_6n152) );
  OAI21_X2 vscale_core_DW01_sub_6_U539 ( .B1(vscale_core_DW01_sub_6n289), .B2(vscale_core_DW01_sub_6n278), .A(vscale_core_DW01_sub_6n279), .ZN(vscale_core_DW01_sub_6n277) );
  OAI21_X2 vscale_core_DW01_sub_6_U540 ( .B1(vscale_core_DW01_sub_6n312), .B2(vscale_core_DW01_sub_6n303), .A(vscale_core_DW01_sub_6n304), .ZN(vscale_core_DW01_sub_6n302) );
  OAI21_X2 vscale_core_DW01_sub_6_U541 ( .B1(vscale_core_DW01_sub_6n174), .B2(vscale_core_DW01_sub_6n124), .A(vscale_core_DW01_sub_6n125), .ZN(vscale_core_DW01_sub_6n123) );
  OAI21_X2 vscale_core_DW01_sub_6_U542 ( .B1(vscale_core_DW01_sub_6n151), .B2(vscale_core_DW01_sub_6n140), .A(vscale_core_DW01_sub_6n141), .ZN(vscale_core_DW01_sub_6n139) );
  OAI21_X2 vscale_core_DW01_sub_6_U543 ( .B1(vscale_core_DW01_sub_6n174), .B2(vscale_core_DW01_sub_6n165), .A(vscale_core_DW01_sub_6n166), .ZN(vscale_core_DW01_sub_6n164) );
  OAI21_X2 vscale_core_DW01_sub_6_U544 ( .B1(vscale_core_DW01_sub_6n174), .B2(vscale_core_DW01_sub_6n112), .A(vscale_core_DW01_sub_6n113), .ZN(vscale_core_DW01_sub_6n111) );
  AOI21_X2 vscale_core_DW01_sub_6_U545 ( .B1(vscale_core_DW01_sub_6n71), .B2(vscale_core_DW01_sub_6n665), .A(vscale_core_DW01_sub_6n68), .ZN(vscale_core_DW01_sub_6n66) );
  AOI21_X2 vscale_core_DW01_sub_6_U546 ( .B1(vscale_core_DW01_sub_6n79), .B2(vscale_core_DW01_sub_6n664), .A(vscale_core_DW01_sub_6n76), .ZN(vscale_core_DW01_sub_6n74) );
  AOI21_X2 vscale_core_DW01_sub_6_U547 ( .B1(vscale_core_DW01_sub_6n87), .B2(vscale_core_DW01_sub_6n662), .A(vscale_core_DW01_sub_6n84), .ZN(vscale_core_DW01_sub_6n82) );
  AOI21_X2 vscale_core_DW01_sub_6_U548 ( .B1(vscale_core_DW01_sub_6n95), .B2(vscale_core_DW01_sub_6n661), .A(vscale_core_DW01_sub_6n92), .ZN(vscale_core_DW01_sub_6n90) );
  AOI21_X2 vscale_core_DW01_sub_6_U549 ( .B1(vscale_core_DW01_sub_6n103), .B2(vscale_core_DW01_sub_6n663), .A(vscale_core_DW01_sub_6n100), .ZN(vscale_core_DW01_sub_6n98) );
  AOI21_X2 vscale_core_DW01_sub_6_U550 ( .B1(vscale_core_DW01_sub_6n175), .B2(vscale_core_DW01_sub_6n107), .A(vscale_core_DW01_sub_6n108), .ZN(vscale_core_DW01_sub_6n106) );
  NOR2_X2 vscale_core_DW01_sub_6_U551 ( .A1(vscale_core_DW01_sub_6n112), .A2(vscale_core_DW01_sub_6n109), .ZN(vscale_core_DW01_sub_6n107) );
  OAI21_X2 vscale_core_DW01_sub_6_U552 ( .B1(vscale_core_DW01_sub_6n113), .B2(vscale_core_DW01_sub_6n109), .A(vscale_core_DW01_sub_6n110), .ZN(vscale_core_DW01_sub_6n108) );
  AOI21_X2 vscale_core_DW01_sub_6_U553 ( .B1(vscale_core_DW01_sub_6n293), .B2(vscale_core_DW01_sub_6n306), .A(vscale_core_DW01_sub_6n294), .ZN(vscale_core_DW01_sub_6n292) );
  OAI21_X2 vscale_core_DW01_sub_6_U554 ( .B1(vscale_core_DW01_sub_6n295), .B2(vscale_core_DW01_sub_6n301), .A(vscale_core_DW01_sub_6n296), .ZN(vscale_core_DW01_sub_6n294) );
  AOI21_X2 vscale_core_DW01_sub_6_U555 ( .B1(vscale_core_DW01_sub_6n155), .B2(vscale_core_DW01_sub_6n168), .A(vscale_core_DW01_sub_6n156), .ZN(vscale_core_DW01_sub_6n154) );
  OAI21_X2 vscale_core_DW01_sub_6_U556 ( .B1(vscale_core_DW01_sub_6n157), .B2(vscale_core_DW01_sub_6n163), .A(vscale_core_DW01_sub_6n158), .ZN(vscale_core_DW01_sub_6n156) );
  AOI21_X2 vscale_core_DW01_sub_6_U557 ( .B1(vscale_core_DW01_sub_6n127), .B2(vscale_core_DW01_sub_6n114), .A(vscale_core_DW01_sub_6n115), .ZN(vscale_core_DW01_sub_6n113) );
  OAI21_X2 vscale_core_DW01_sub_6_U558 ( .B1(vscale_core_DW01_sub_6n116), .B2(vscale_core_DW01_sub_6n122), .A(vscale_core_DW01_sub_6n117), .ZN(vscale_core_DW01_sub_6n115) );
  AOI21_X2 vscale_core_DW01_sub_6_U559 ( .B1(vscale_core_DW01_sub_6n203), .B2(vscale_core_DW01_sub_6n212), .A(vscale_core_DW01_sub_6n204), .ZN(vscale_core_DW01_sub_6n202) );
  OAI21_X2 vscale_core_DW01_sub_6_U560 ( .B1(vscale_core_DW01_sub_6n205), .B2(vscale_core_DW01_sub_6n209), .A(vscale_core_DW01_sub_6n206), .ZN(vscale_core_DW01_sub_6n204) );
  AOI21_X2 vscale_core_DW01_sub_6_U561 ( .B1(vscale_core_DW01_sub_6n245), .B2(vscale_core_DW01_sub_6n254), .A(vscale_core_DW01_sub_6n246), .ZN(vscale_core_DW01_sub_6n244) );
  OAI21_X2 vscale_core_DW01_sub_6_U562 ( .B1(vscale_core_DW01_sub_6n247), .B2(vscale_core_DW01_sub_6n251), .A(vscale_core_DW01_sub_6n248), .ZN(vscale_core_DW01_sub_6n246) );
  OAI21_X2 vscale_core_DW01_sub_6_U563 ( .B1(vscale_core_DW01_sub_6n244), .B2(vscale_core_DW01_sub_6n222), .A(vscale_core_DW01_sub_6n223), .ZN(vscale_core_DW01_sub_6n221) );
  AOI21_X2 vscale_core_DW01_sub_6_U564 ( .B1(vscale_core_DW01_sub_6n224), .B2(vscale_core_DW01_sub_6n233), .A(vscale_core_DW01_sub_6n225), .ZN(vscale_core_DW01_sub_6n223) );
  OAI21_X2 vscale_core_DW01_sub_6_U565 ( .B1(vscale_core_DW01_sub_6n226), .B2(vscale_core_DW01_sub_6n230), .A(vscale_core_DW01_sub_6n227), .ZN(vscale_core_DW01_sub_6n225) );
  OAI21_X2 vscale_core_DW01_sub_6_U566 ( .B1(vscale_core_DW01_sub_6n334), .B2(vscale_core_DW01_sub_6n314), .A(vscale_core_DW01_sub_6n315), .ZN(vscale_core_DW01_sub_6n313) );
  AOI21_X2 vscale_core_DW01_sub_6_U567 ( .B1(vscale_core_DW01_sub_6n316), .B2(vscale_core_DW01_sub_6n325), .A(vscale_core_DW01_sub_6n317), .ZN(vscale_core_DW01_sub_6n315) );
  NOR2_X2 vscale_core_DW01_sub_6_U568 ( .A1(vscale_core_DW01_sub_6n318), .A2(vscale_core_DW01_sub_6n321), .ZN(vscale_core_DW01_sub_6n316) );
  OAI21_X2 vscale_core_DW01_sub_6_U569 ( .B1(vscale_core_DW01_sub_6n154), .B2(vscale_core_DW01_sub_6n128), .A(vscale_core_DW01_sub_6n129), .ZN(vscale_core_DW01_sub_6n127) );
  AOI21_X2 vscale_core_DW01_sub_6_U570 ( .B1(vscale_core_DW01_sub_6n130), .B2(vscale_core_DW01_sub_6n143), .A(vscale_core_DW01_sub_6n131), .ZN(vscale_core_DW01_sub_6n129) );
  OAI21_X2 vscale_core_DW01_sub_6_U571 ( .B1(vscale_core_DW01_sub_6n132), .B2(vscale_core_DW01_sub_6n138), .A(vscale_core_DW01_sub_6n133), .ZN(vscale_core_DW01_sub_6n131) );
  OAI21_X2 vscale_core_DW01_sub_6_U572 ( .B1(vscale_core_DW01_sub_6n74), .B2(vscale_core_DW01_sub_6n72), .A(vscale_core_DW01_sub_6n73), .ZN(vscale_core_DW01_sub_6n71) );
  OAI21_X2 vscale_core_DW01_sub_6_U573 ( .B1(vscale_core_DW01_sub_6n82), .B2(vscale_core_DW01_sub_6n80), .A(vscale_core_DW01_sub_6n81), .ZN(vscale_core_DW01_sub_6n79) );
  OAI21_X2 vscale_core_DW01_sub_6_U574 ( .B1(vscale_core_DW01_sub_6n90), .B2(vscale_core_DW01_sub_6n88), .A(vscale_core_DW01_sub_6n89), .ZN(vscale_core_DW01_sub_6n87) );
  OAI21_X2 vscale_core_DW01_sub_6_U575 ( .B1(vscale_core_DW01_sub_6n98), .B2(vscale_core_DW01_sub_6n96), .A(vscale_core_DW01_sub_6n97), .ZN(vscale_core_DW01_sub_6n95) );
  OAI21_X2 vscale_core_DW01_sub_6_U576 ( .B1(vscale_core_DW01_sub_6n106), .B2(vscale_core_DW01_sub_6n104), .A(vscale_core_DW01_sub_6n105), .ZN(vscale_core_DW01_sub_6n103) );
  OAI21_X2 vscale_core_DW01_sub_6_U577 ( .B1(vscale_core_DW01_sub_6n326), .B2(vscale_core_DW01_sub_6n332), .A(vscale_core_DW01_sub_6n327), .ZN(vscale_core_DW01_sub_6n325) );
  OAI21_X2 vscale_core_DW01_sub_6_U578 ( .B1(vscale_core_DW01_sub_6n213), .B2(vscale_core_DW01_sub_6n217), .A(vscale_core_DW01_sub_6n214), .ZN(vscale_core_DW01_sub_6n212) );
  OAI21_X2 vscale_core_DW01_sub_6_U579 ( .B1(vscale_core_DW01_sub_6n255), .B2(vscale_core_DW01_sub_6n261), .A(vscale_core_DW01_sub_6n256), .ZN(vscale_core_DW01_sub_6n254) );
  OAI21_X2 vscale_core_DW01_sub_6_U580 ( .B1(vscale_core_DW01_sub_6n192), .B2(vscale_core_DW01_sub_6n196), .A(vscale_core_DW01_sub_6n193), .ZN(vscale_core_DW01_sub_6n191) );
  OAI21_X2 vscale_core_DW01_sub_6_U581 ( .B1(vscale_core_DW01_sub_6n234), .B2(vscale_core_DW01_sub_6n238), .A(vscale_core_DW01_sub_6n235), .ZN(vscale_core_DW01_sub_6n233) );
  OAI21_X2 vscale_core_DW01_sub_6_U582 ( .B1(vscale_core_DW01_sub_6n307), .B2(vscale_core_DW01_sub_6n311), .A(vscale_core_DW01_sub_6n308), .ZN(vscale_core_DW01_sub_6n306) );
  OAI21_X2 vscale_core_DW01_sub_6_U583 ( .B1(vscale_core_DW01_sub_6n282), .B2(vscale_core_DW01_sub_6n288), .A(vscale_core_DW01_sub_6n283), .ZN(vscale_core_DW01_sub_6n281) );
  OAI21_X2 vscale_core_DW01_sub_6_U584 ( .B1(vscale_core_DW01_sub_6n344), .B2(vscale_core_DW01_sub_6n346), .A(vscale_core_DW01_sub_6n345), .ZN(vscale_core_DW01_sub_6n343) );
  OAI21_X2 vscale_core_DW01_sub_6_U585 ( .B1(vscale_core_DW01_sub_6n169), .B2(vscale_core_DW01_sub_6n173), .A(vscale_core_DW01_sub_6n170), .ZN(vscale_core_DW01_sub_6n168) );
  OAI21_X2 vscale_core_DW01_sub_6_U586 ( .B1(vscale_core_DW01_sub_6n144), .B2(vscale_core_DW01_sub_6n150), .A(vscale_core_DW01_sub_6n145), .ZN(vscale_core_DW01_sub_6n143) );
  AOI21_X2 vscale_core_DW01_sub_6_U587 ( .B1(vscale_core_DW01_sub_6n268), .B2(vscale_core_DW01_sub_6n281), .A(vscale_core_DW01_sub_6n269), .ZN(vscale_core_DW01_sub_6n267) );
  OAI21_X2 vscale_core_DW01_sub_6_U588 ( .B1(vscale_core_DW01_sub_6n270), .B2(vscale_core_DW01_sub_6n276), .A(vscale_core_DW01_sub_6n271), .ZN(vscale_core_DW01_sub_6n269) );
  OAI21_X2 vscale_core_DW01_sub_6_U589 ( .B1(vscale_core_DW01_sub_6n318), .B2(vscale_core_DW01_sub_6n322), .A(vscale_core_DW01_sub_6n319), .ZN(vscale_core_DW01_sub_6n317) );
  AOI21_X2 vscale_core_DW01_sub_6_U590 ( .B1(vscale_core_DW01_sub_6n335), .B2(vscale_core_DW01_sub_6n343), .A(vscale_core_DW01_sub_6n336), .ZN(vscale_core_DW01_sub_6n334) );
  NOR2_X2 vscale_core_DW01_sub_6_U591 ( .A1(vscale_core_DW01_sub_6n337), .A2(vscale_core_DW01_sub_6n340), .ZN(vscale_core_DW01_sub_6n335) );
  OAI21_X2 vscale_core_DW01_sub_6_U592 ( .B1(vscale_core_DW01_sub_6n337), .B2(vscale_core_DW01_sub_6n341), .A(vscale_core_DW01_sub_6n338), .ZN(vscale_core_DW01_sub_6n336) );
  OAI21_X2 vscale_core_DW01_sub_6_U593 ( .B1(vscale_core_DW01_sub_6n202), .B2(vscale_core_DW01_sub_6n180), .A(vscale_core_DW01_sub_6n181), .ZN(vscale_core_DW01_sub_6n179) );
  AOI21_X2 vscale_core_DW01_sub_6_U594 ( .B1(vscale_core_DW01_sub_6n182), .B2(vscale_core_DW01_sub_6n191), .A(vscale_core_DW01_sub_6n183), .ZN(vscale_core_DW01_sub_6n181) );
  OAI21_X2 vscale_core_DW01_sub_6_U595 ( .B1(vscale_core_DW01_sub_6n184), .B2(vscale_core_DW01_sub_6n188), .A(vscale_core_DW01_sub_6n185), .ZN(vscale_core_DW01_sub_6n183) );
  NOR2_X2 vscale_core_DW01_sub_6_U596 ( .A1(vscale_core_DW01_sub_6n270), .A2(vscale_core_DW01_sub_6n275), .ZN(vscale_core_DW01_sub_6n268) );
  NOR2_X2 vscale_core_DW01_sub_6_U597 ( .A1(vscale_core_DW01_sub_6n295), .A2(vscale_core_DW01_sub_6n300), .ZN(vscale_core_DW01_sub_6n293) );
  NOR2_X2 vscale_core_DW01_sub_6_U598 ( .A1(vscale_core_DW01_sub_6n205), .A2(vscale_core_DW01_sub_6n208), .ZN(vscale_core_DW01_sub_6n203) );
  NOR2_X2 vscale_core_DW01_sub_6_U599 ( .A1(vscale_core_DW01_sub_6n226), .A2(vscale_core_DW01_sub_6n229), .ZN(vscale_core_DW01_sub_6n224) );
  NOR2_X2 vscale_core_DW01_sub_6_U600 ( .A1(vscale_core_DW01_sub_6n247), .A2(vscale_core_DW01_sub_6n250), .ZN(vscale_core_DW01_sub_6n245) );
  NOR2_X2 vscale_core_DW01_sub_6_U601 ( .A1(vscale_core_DW01_sub_6n132), .A2(vscale_core_DW01_sub_6n137), .ZN(vscale_core_DW01_sub_6n130) );
  NOR2_X2 vscale_core_DW01_sub_6_U602 ( .A1(vscale_core_DW01_sub_6n157), .A2(vscale_core_DW01_sub_6n162), .ZN(vscale_core_DW01_sub_6n155) );
  NOR2_X2 vscale_core_DW01_sub_6_U603 ( .A1(vscale_core_DW01_sub_6n184), .A2(vscale_core_DW01_sub_6n187), .ZN(vscale_core_DW01_sub_6n182) );
  NOR2_X2 vscale_core_DW01_sub_6_U604 ( .A1(vscale_core_DW01_sub_6n192), .A2(vscale_core_DW01_sub_6n195), .ZN(vscale_core_DW01_sub_6n190) );
  NOR2_X2 vscale_core_DW01_sub_6_U605 ( .A1(vscale_core_DW01_sub_6n282), .A2(vscale_core_DW01_sub_6n287), .ZN(vscale_core_DW01_sub_6n280) );
  NOR2_X2 vscale_core_DW01_sub_6_U606 ( .A1(vscale_core_DW01_sub_6n144), .A2(vscale_core_DW01_sub_6n149), .ZN(vscale_core_DW01_sub_6n142) );
  NOR2_X2 vscale_core_DW01_sub_6_U607 ( .A1(vscale_core_DW01_sub_6n331), .A2(vscale_core_DW01_sub_6n326), .ZN(vscale_core_DW01_sub_6n324) );
  NOR2_X2 vscale_core_DW01_sub_6_U608 ( .A1(vscale_core_DW01_sub_6n234), .A2(vscale_core_DW01_sub_6n237), .ZN(vscale_core_DW01_sub_6n232) );
  NOR2_X2 vscale_core_DW01_sub_6_U609 ( .A1(vscale_core_DW01_sub_6n255), .A2(vscale_core_DW01_sub_6n260), .ZN(vscale_core_DW01_sub_6n253) );
  NOR2_X2 vscale_core_DW01_sub_6_U610 ( .A1(vscale_core_DW01_sub_6n213), .A2(vscale_core_DW01_sub_6n216), .ZN(vscale_core_DW01_sub_6n211) );
  NOR2_X2 vscale_core_DW01_sub_6_U611 ( .A1(vscale_core_DW01_sub_6n116), .A2(vscale_core_DW01_sub_6n121), .ZN(vscale_core_DW01_sub_6n114) );
  NOR2_X2 vscale_core_DW01_sub_6_U612 ( .A1(vscale_core_DW01_sub_6n307), .A2(vscale_core_DW01_sub_6n310), .ZN(vscale_core_DW01_sub_6n305) );
  NOR2_X2 vscale_core_DW01_sub_6_U613 ( .A1(vscale_core_DW01_sub_6n169), .A2(vscale_core_DW01_sub_6n172), .ZN(vscale_core_DW01_sub_6n167) );
  OAI21_X2 vscale_core_DW01_sub_6_U614 ( .B1(vscale_core_DW01_sub_6n189), .B2(vscale_core_DW01_sub_6n187), .A(vscale_core_DW01_sub_6n188), .ZN(vscale_core_DW01_sub_6n186) );
  AOI21_X2 vscale_core_DW01_sub_6_U615 ( .B1(vscale_core_DW01_sub_6n262), .B2(vscale_core_DW01_sub_6n384), .A(vscale_core_DW01_sub_6n259), .ZN(vscale_core_DW01_sub_6n257) );
  AOI21_X2 vscale_core_DW01_sub_6_U616 ( .B1(vscale_core_DW01_sub_6n277), .B2(vscale_core_DW01_sub_6n386), .A(vscale_core_DW01_sub_6n274), .ZN(vscale_core_DW01_sub_6n272) );
  AOI21_X2 vscale_core_DW01_sub_6_U617 ( .B1(vscale_core_DW01_sub_6n290), .B2(vscale_core_DW01_sub_6n388), .A(vscale_core_DW01_sub_6n286), .ZN(vscale_core_DW01_sub_6n284) );
  AOI21_X2 vscale_core_DW01_sub_6_U618 ( .B1(vscale_core_DW01_sub_6n302), .B2(vscale_core_DW01_sub_6n390), .A(vscale_core_DW01_sub_6n299), .ZN(vscale_core_DW01_sub_6n297) );
  AOI21_X2 vscale_core_DW01_sub_6_U619 ( .B1(vscale_core_DW01_sub_6n123), .B2(vscale_core_DW01_sub_6n360), .A(vscale_core_DW01_sub_6n120), .ZN(vscale_core_DW01_sub_6n118) );
  AOI21_X2 vscale_core_DW01_sub_6_U620 ( .B1(vscale_core_DW01_sub_6n139), .B2(vscale_core_DW01_sub_6n362), .A(vscale_core_DW01_sub_6n136), .ZN(vscale_core_DW01_sub_6n134) );
  AOI21_X2 vscale_core_DW01_sub_6_U621 ( .B1(vscale_core_DW01_sub_6n152), .B2(vscale_core_DW01_sub_6n364), .A(vscale_core_DW01_sub_6n148), .ZN(vscale_core_DW01_sub_6n146) );
  AOI21_X2 vscale_core_DW01_sub_6_U622 ( .B1(vscale_core_DW01_sub_6n164), .B2(vscale_core_DW01_sub_6n366), .A(vscale_core_DW01_sub_6n161), .ZN(vscale_core_DW01_sub_6n159) );
  OAI21_X2 vscale_core_DW01_sub_6_U623 ( .B1(vscale_core_DW01_sub_6n198), .B2(vscale_core_DW01_sub_6n195), .A(vscale_core_DW01_sub_6n196), .ZN(vscale_core_DW01_sub_6n194) );
  OAI21_X2 vscale_core_DW01_sub_6_U624 ( .B1(vscale_core_DW01_sub_6n210), .B2(vscale_core_DW01_sub_6n208), .A(vscale_core_DW01_sub_6n209), .ZN(vscale_core_DW01_sub_6n207) );
  OAI21_X2 vscale_core_DW01_sub_6_U625 ( .B1(vscale_core_DW01_sub_6n219), .B2(vscale_core_DW01_sub_6n216), .A(vscale_core_DW01_sub_6n217), .ZN(vscale_core_DW01_sub_6n215) );
  OAI21_X2 vscale_core_DW01_sub_6_U626 ( .B1(vscale_core_DW01_sub_6n231), .B2(vscale_core_DW01_sub_6n229), .A(vscale_core_DW01_sub_6n230), .ZN(vscale_core_DW01_sub_6n228) );
  OAI21_X2 vscale_core_DW01_sub_6_U627 ( .B1(vscale_core_DW01_sub_6n240), .B2(vscale_core_DW01_sub_6n237), .A(vscale_core_DW01_sub_6n238), .ZN(vscale_core_DW01_sub_6n236) );
  OAI21_X2 vscale_core_DW01_sub_6_U628 ( .B1(vscale_core_DW01_sub_6n252), .B2(vscale_core_DW01_sub_6n250), .A(vscale_core_DW01_sub_6n251), .ZN(vscale_core_DW01_sub_6n249) );
  OAI21_X2 vscale_core_DW01_sub_6_U629 ( .B1(vscale_core_DW01_sub_6n312), .B2(vscale_core_DW01_sub_6n310), .A(vscale_core_DW01_sub_6n311), .ZN(vscale_core_DW01_sub_6n309) );
  OAI21_X2 vscale_core_DW01_sub_6_U630 ( .B1(vscale_core_DW01_sub_6n323), .B2(vscale_core_DW01_sub_6n321), .A(vscale_core_DW01_sub_6n322), .ZN(vscale_core_DW01_sub_6n320) );
  AOI21_X2 vscale_core_DW01_sub_6_U631 ( .B1(vscale_core_DW01_sub_6n333), .B2(vscale_core_DW01_sub_6n396), .A(vscale_core_DW01_sub_6n330), .ZN(vscale_core_DW01_sub_6n328) );
  OAI21_X2 vscale_core_DW01_sub_6_U632 ( .B1(vscale_core_DW01_sub_6n342), .B2(vscale_core_DW01_sub_6n340), .A(vscale_core_DW01_sub_6n341), .ZN(vscale_core_DW01_sub_6n339) );
  OAI21_X2 vscale_core_DW01_sub_6_U633 ( .B1(vscale_core_DW01_sub_6n174), .B2(vscale_core_DW01_sub_6n172), .A(vscale_core_DW01_sub_6n173), .ZN(vscale_core_DW01_sub_6n171) );
  NOR2_X2 vscale_core_DW01_sub_6_U634 ( .A1(vscale_core_DW01_sub_6n459), .A2(pipeline_md_a[3]), .ZN(vscale_core_DW01_sub_6n337) );
  NOR2_X2 vscale_core_DW01_sub_6_U635 ( .A1(vscale_core_DW01_sub_6n455), .A2(pipeline_md_a[7]), .ZN(vscale_core_DW01_sub_6n318) );
  NOR2_X2 vscale_core_DW01_sub_6_U636 ( .A1(vscale_core_DW01_sub_6n447), .A2(pipeline_md_a[15]), .ZN(vscale_core_DW01_sub_6n270) );
  NOR2_X2 vscale_core_DW01_sub_6_U637 ( .A1(vscale_core_DW01_sub_6n449), .A2(pipeline_md_a[13]), .ZN(vscale_core_DW01_sub_6n282) );
  NOR2_X2 vscale_core_DW01_sub_6_U638 ( .A1(vscale_core_DW01_sub_6n451), .A2(pipeline_md_a[11]), .ZN(vscale_core_DW01_sub_6n295) );
  NOR2_X2 vscale_core_DW01_sub_6_U639 ( .A1(vscale_core_DW01_sub_6n453), .A2(pipeline_md_a[9]), .ZN(vscale_core_DW01_sub_6n307) );
  NOR2_X2 vscale_core_DW01_sub_6_U640 ( .A1(vscale_core_DW01_sub_6n423), .A2(pipeline_md_a[39]), .ZN(vscale_core_DW01_sub_6n132) );
  NOR2_X2 vscale_core_DW01_sub_6_U641 ( .A1(vscale_core_DW01_sub_6n425), .A2(pipeline_md_a[37]), .ZN(vscale_core_DW01_sub_6n144) );
  NOR2_X2 vscale_core_DW01_sub_6_U642 ( .A1(vscale_core_DW01_sub_6n427), .A2(pipeline_md_a[35]), .ZN(vscale_core_DW01_sub_6n157) );
  NOR2_X2 vscale_core_DW01_sub_6_U643 ( .A1(vscale_core_DW01_sub_6n429), .A2(pipeline_md_a[33]), .ZN(vscale_core_DW01_sub_6n169) );
  NOR2_X2 vscale_core_DW01_sub_6_U644 ( .A1(vscale_core_DW01_sub_6n431), .A2(pipeline_md_a[31]), .ZN(vscale_core_DW01_sub_6n184) );
  NOR2_X2 vscale_core_DW01_sub_6_U645 ( .A1(vscale_core_DW01_sub_6n433), .A2(pipeline_md_a[29]), .ZN(vscale_core_DW01_sub_6n192) );
  NOR2_X2 vscale_core_DW01_sub_6_U646 ( .A1(vscale_core_DW01_sub_6n435), .A2(pipeline_md_a[27]), .ZN(vscale_core_DW01_sub_6n205) );
  NOR2_X2 vscale_core_DW01_sub_6_U647 ( .A1(vscale_core_DW01_sub_6n437), .A2(pipeline_md_a[25]), .ZN(vscale_core_DW01_sub_6n213) );
  NOR2_X2 vscale_core_DW01_sub_6_U648 ( .A1(vscale_core_DW01_sub_6n439), .A2(pipeline_md_a[23]), .ZN(vscale_core_DW01_sub_6n226) );
  NOR2_X2 vscale_core_DW01_sub_6_U649 ( .A1(vscale_core_DW01_sub_6n441), .A2(pipeline_md_a[21]), .ZN(vscale_core_DW01_sub_6n234) );
  NOR2_X2 vscale_core_DW01_sub_6_U650 ( .A1(vscale_core_DW01_sub_6n443), .A2(pipeline_md_a[19]), .ZN(vscale_core_DW01_sub_6n247) );
  NOR2_X2 vscale_core_DW01_sub_6_U651 ( .A1(vscale_core_DW01_sub_6n445), .A2(pipeline_md_a[17]), .ZN(vscale_core_DW01_sub_6n255) );
  NOR2_X2 vscale_core_DW01_sub_6_U652 ( .A1(vscale_core_DW01_sub_6n457), .A2(pipeline_md_a[5]), .ZN(vscale_core_DW01_sub_6n326) );
  OAI21_X2 vscale_core_DW01_sub_6_U653 ( .B1(vscale_core_DW01_sub_6n66), .B2(vscale_core_DW01_sub_6n64), .A(vscale_core_DW01_sub_6n65), .ZN(vscale_core_DW01_sub_6n63) );
  NOR2_X2 vscale_core_DW01_sub_6_U654 ( .A1(vscale_core_DW01_sub_6n434), .A2(pipeline_md_a[28]), .ZN(vscale_core_DW01_sub_6n195) );
  NOR2_X2 vscale_core_DW01_sub_6_U655 ( .A1(vscale_core_DW01_sub_6n436), .A2(pipeline_md_a[26]), .ZN(vscale_core_DW01_sub_6n208) );
  NOR2_X2 vscale_core_DW01_sub_6_U656 ( .A1(vscale_core_DW01_sub_6n440), .A2(pipeline_md_a[22]), .ZN(vscale_core_DW01_sub_6n229) );
  NOR2_X2 vscale_core_DW01_sub_6_U657 ( .A1(vscale_core_DW01_sub_6n444), .A2(pipeline_md_a[18]), .ZN(vscale_core_DW01_sub_6n250) );
  NOR2_X2 vscale_core_DW01_sub_6_U658 ( .A1(vscale_core_DW01_sub_6n456), .A2(pipeline_md_a[6]), .ZN(vscale_core_DW01_sub_6n321) );
  NOR2_X2 vscale_core_DW01_sub_6_U659 ( .A1(vscale_core_DW01_sub_6n460), .A2(pipeline_md_a[2]), .ZN(vscale_core_DW01_sub_6n340) );
  NOR2_X2 vscale_core_DW01_sub_6_U660 ( .A1(vscale_core_DW01_sub_6n432), .A2(pipeline_md_a[30]), .ZN(vscale_core_DW01_sub_6n187) );
  NOR2_X2 vscale_core_DW01_sub_6_U661 ( .A1(vscale_core_DW01_sub_6n461), .A2(pipeline_md_a[1]), .ZN(vscale_core_DW01_sub_6n344) );
  NOR2_X2 vscale_core_DW01_sub_6_U662 ( .A1(vscale_core_DW01_sub_6n448), .A2(pipeline_md_a[14]), .ZN(vscale_core_DW01_sub_6n275) );
  NOR2_X2 vscale_core_DW01_sub_6_U663 ( .A1(vscale_core_DW01_sub_6n450), .A2(pipeline_md_a[12]), .ZN(vscale_core_DW01_sub_6n287) );
  NOR2_X2 vscale_core_DW01_sub_6_U664 ( .A1(vscale_core_DW01_sub_6n452), .A2(pipeline_md_a[10]), .ZN(vscale_core_DW01_sub_6n300) );
  NOR2_X2 vscale_core_DW01_sub_6_U665 ( .A1(vscale_core_DW01_sub_6n424), .A2(pipeline_md_a[38]), .ZN(vscale_core_DW01_sub_6n137) );
  NOR2_X2 vscale_core_DW01_sub_6_U666 ( .A1(vscale_core_DW01_sub_6n426), .A2(pipeline_md_a[36]), .ZN(vscale_core_DW01_sub_6n149) );
  NOR2_X2 vscale_core_DW01_sub_6_U667 ( .A1(vscale_core_DW01_sub_6n428), .A2(pipeline_md_a[34]), .ZN(vscale_core_DW01_sub_6n162) );
  NOR2_X2 vscale_core_DW01_sub_6_U668 ( .A1(vscale_core_DW01_sub_6n462), .A2(pipeline_md_a[0]), .ZN(vscale_core_DW01_sub_6n346) );
  NOR2_X2 vscale_core_DW01_sub_6_U669 ( .A1(vscale_core_DW01_sub_6n421), .A2(pipeline_md_a[41]), .ZN(vscale_core_DW01_sub_6n116) );
  NOR2_X2 vscale_core_DW01_sub_6_U670 ( .A1(vscale_core_DW01_sub_6n438), .A2(pipeline_md_a[24]), .ZN(vscale_core_DW01_sub_6n216) );
  NOR2_X2 vscale_core_DW01_sub_6_U671 ( .A1(vscale_core_DW01_sub_6n442), .A2(pipeline_md_a[20]), .ZN(vscale_core_DW01_sub_6n237) );
  NOR2_X2 vscale_core_DW01_sub_6_U672 ( .A1(vscale_core_DW01_sub_6n454), .A2(pipeline_md_a[8]), .ZN(vscale_core_DW01_sub_6n310) );
  NOR2_X2 vscale_core_DW01_sub_6_U673 ( .A1(vscale_core_DW01_sub_6n420), .A2(pipeline_md_a[42]), .ZN(vscale_core_DW01_sub_6n109) );
  NOR2_X2 vscale_core_DW01_sub_6_U674 ( .A1(vscale_core_DW01_sub_6n430), .A2(pipeline_md_a[32]), .ZN(vscale_core_DW01_sub_6n172) );
  NOR2_X2 vscale_core_DW01_sub_6_U675 ( .A1(vscale_core_DW01_sub_6n458), .A2(pipeline_md_a[4]), .ZN(vscale_core_DW01_sub_6n331) );
  NOR2_X2 vscale_core_DW01_sub_6_U676 ( .A1(vscale_core_DW01_sub_6n446), .A2(pipeline_md_a[16]), .ZN(vscale_core_DW01_sub_6n260) );
  NOR2_X2 vscale_core_DW01_sub_6_U677 ( .A1(vscale_core_DW01_sub_6n422), .A2(pipeline_md_a[40]), .ZN(vscale_core_DW01_sub_6n121) );
  NOR2_X2 vscale_core_DW01_sub_6_U678 ( .A1(vscale_core_DW01_sub_6n419), .A2(pipeline_md_a[43]), .ZN(vscale_core_DW01_sub_6n104) );
  NOR2_X2 vscale_core_DW01_sub_6_U679 ( .A1(vscale_core_DW01_sub_6n413), .A2(pipeline_md_a[49]), .ZN(vscale_core_DW01_sub_6n80) );
  NOR2_X2 vscale_core_DW01_sub_6_U680 ( .A1(vscale_core_DW01_sub_6n415), .A2(pipeline_md_a[47]), .ZN(vscale_core_DW01_sub_6n88) );
  NOR2_X2 vscale_core_DW01_sub_6_U681 ( .A1(vscale_core_DW01_sub_6n417), .A2(pipeline_md_a[45]), .ZN(vscale_core_DW01_sub_6n96) );
  OR2_X1 vscale_core_DW01_sub_6_U682 ( .A1(vscale_core_DW01_sub_6n416), .A2(pipeline_md_a[46]), .ZN(vscale_core_DW01_sub_6n661) );
  OR2_X1 vscale_core_DW01_sub_6_U683 ( .A1(vscale_core_DW01_sub_6n414), .A2(pipeline_md_a[48]), .ZN(vscale_core_DW01_sub_6n662) );
  OR2_X1 vscale_core_DW01_sub_6_U684 ( .A1(vscale_core_DW01_sub_6n418), .A2(pipeline_md_a[44]), .ZN(vscale_core_DW01_sub_6n663) );
  NOR2_X2 vscale_core_DW01_sub_6_U685 ( .A1(vscale_core_DW01_sub_6n409), .A2(pipeline_md_a[53]), .ZN(vscale_core_DW01_sub_6n64) );
  NOR2_X2 vscale_core_DW01_sub_6_U686 ( .A1(vscale_core_DW01_sub_6n411), .A2(pipeline_md_a[51]), .ZN(vscale_core_DW01_sub_6n72) );
  OR2_X1 vscale_core_DW01_sub_6_U687 ( .A1(vscale_core_DW01_sub_6n412), .A2(pipeline_md_a[50]), .ZN(vscale_core_DW01_sub_6n664) );
  OR2_X1 vscale_core_DW01_sub_6_U688 ( .A1(vscale_core_DW01_sub_6n410), .A2(pipeline_md_a[52]), .ZN(vscale_core_DW01_sub_6n665) );
  INV_X4 vscale_core_DW01_sub_6_U689 ( .A(vscale_core_DW01_sub_6n94), .ZN(vscale_core_DW01_sub_6n92) );
  INV_X4 vscale_core_DW01_sub_6_U690 ( .A(vscale_core_DW01_sub_6n86), .ZN(vscale_core_DW01_sub_6n84) );
  INV_X4 vscale_core_DW01_sub_6_U691 ( .A(vscale_core_DW01_sub_6n78), .ZN(vscale_core_DW01_sub_6n76) );
  INV_X4 vscale_core_DW01_sub_6_U692 ( .A(vscale_core_DW01_sub_6n70), .ZN(vscale_core_DW01_sub_6n68) );
  INV_X4 vscale_core_DW01_sub_6_U693 ( .A(pipeline_md_b[0]), .ZN(vscale_core_DW01_sub_6n462) );
  INV_X4 vscale_core_DW01_sub_6_U694 ( .A(pipeline_md_b[1]), .ZN(vscale_core_DW01_sub_6n461) );
  INV_X4 vscale_core_DW01_sub_6_U695 ( .A(pipeline_md_b[2]), .ZN(vscale_core_DW01_sub_6n460) );
  INV_X4 vscale_core_DW01_sub_6_U696 ( .A(pipeline_md_b[3]), .ZN(vscale_core_DW01_sub_6n459) );
  INV_X4 vscale_core_DW01_sub_6_U697 ( .A(pipeline_md_b[4]), .ZN(vscale_core_DW01_sub_6n458) );
  INV_X4 vscale_core_DW01_sub_6_U698 ( .A(pipeline_md_b[5]), .ZN(vscale_core_DW01_sub_6n457) );
  INV_X4 vscale_core_DW01_sub_6_U699 ( .A(pipeline_md_b[6]), .ZN(vscale_core_DW01_sub_6n456) );
  INV_X4 vscale_core_DW01_sub_6_U700 ( .A(pipeline_md_b[7]), .ZN(vscale_core_DW01_sub_6n455) );
  INV_X4 vscale_core_DW01_sub_6_U701 ( .A(pipeline_md_b[8]), .ZN(vscale_core_DW01_sub_6n454) );
  INV_X4 vscale_core_DW01_sub_6_U702 ( .A(pipeline_md_b[9]), .ZN(vscale_core_DW01_sub_6n453) );
  INV_X4 vscale_core_DW01_sub_6_U703 ( .A(pipeline_md_b[10]), .ZN(vscale_core_DW01_sub_6n452) );
  INV_X4 vscale_core_DW01_sub_6_U704 ( .A(pipeline_md_b[11]), .ZN(vscale_core_DW01_sub_6n451) );
  INV_X4 vscale_core_DW01_sub_6_U705 ( .A(pipeline_md_b[12]), .ZN(vscale_core_DW01_sub_6n450) );
  INV_X4 vscale_core_DW01_sub_6_U706 ( .A(pipeline_md_b[13]), .ZN(vscale_core_DW01_sub_6n449) );
  INV_X4 vscale_core_DW01_sub_6_U707 ( .A(pipeline_md_b[14]), .ZN(vscale_core_DW01_sub_6n448) );
  INV_X4 vscale_core_DW01_sub_6_U708 ( .A(pipeline_md_b[15]), .ZN(vscale_core_DW01_sub_6n447) );
  INV_X4 vscale_core_DW01_sub_6_U709 ( .A(pipeline_md_b[16]), .ZN(vscale_core_DW01_sub_6n446) );
  INV_X4 vscale_core_DW01_sub_6_U710 ( .A(pipeline_md_b[17]), .ZN(vscale_core_DW01_sub_6n445) );
  INV_X4 vscale_core_DW01_sub_6_U711 ( .A(pipeline_md_b[18]), .ZN(vscale_core_DW01_sub_6n444) );
  INV_X4 vscale_core_DW01_sub_6_U712 ( .A(pipeline_md_b[19]), .ZN(vscale_core_DW01_sub_6n443) );
  INV_X4 vscale_core_DW01_sub_6_U713 ( .A(pipeline_md_b[20]), .ZN(vscale_core_DW01_sub_6n442) );
  INV_X4 vscale_core_DW01_sub_6_U714 ( .A(pipeline_md_b[21]), .ZN(vscale_core_DW01_sub_6n441) );
  INV_X4 vscale_core_DW01_sub_6_U715 ( .A(pipeline_md_b[22]), .ZN(vscale_core_DW01_sub_6n440) );
  INV_X4 vscale_core_DW01_sub_6_U716 ( .A(pipeline_md_b[23]), .ZN(vscale_core_DW01_sub_6n439) );
  INV_X4 vscale_core_DW01_sub_6_U717 ( .A(pipeline_md_b[24]), .ZN(vscale_core_DW01_sub_6n438) );
  INV_X4 vscale_core_DW01_sub_6_U718 ( .A(pipeline_md_b[25]), .ZN(vscale_core_DW01_sub_6n437) );
  INV_X4 vscale_core_DW01_sub_6_U719 ( .A(pipeline_md_b[26]), .ZN(vscale_core_DW01_sub_6n436) );
  INV_X4 vscale_core_DW01_sub_6_U720 ( .A(pipeline_md_b[27]), .ZN(vscale_core_DW01_sub_6n435) );
  INV_X4 vscale_core_DW01_sub_6_U721 ( .A(pipeline_md_b[28]), .ZN(vscale_core_DW01_sub_6n434) );
  INV_X4 vscale_core_DW01_sub_6_U722 ( .A(pipeline_md_b[29]), .ZN(vscale_core_DW01_sub_6n433) );
  INV_X4 vscale_core_DW01_sub_6_U723 ( .A(pipeline_md_b[30]), .ZN(vscale_core_DW01_sub_6n432) );
  INV_X4 vscale_core_DW01_sub_6_U724 ( .A(pipeline_md_b[31]), .ZN(vscale_core_DW01_sub_6n431) );
  INV_X4 vscale_core_DW01_sub_6_U725 ( .A(pipeline_md_b[32]), .ZN(vscale_core_DW01_sub_6n430) );
  INV_X4 vscale_core_DW01_sub_6_U726 ( .A(pipeline_md_b[33]), .ZN(vscale_core_DW01_sub_6n429) );
  INV_X4 vscale_core_DW01_sub_6_U727 ( .A(pipeline_md_b[34]), .ZN(vscale_core_DW01_sub_6n428) );
  INV_X4 vscale_core_DW01_sub_6_U728 ( .A(pipeline_md_b[35]), .ZN(vscale_core_DW01_sub_6n427) );
  INV_X4 vscale_core_DW01_sub_6_U729 ( .A(pipeline_md_b[36]), .ZN(vscale_core_DW01_sub_6n426) );
  INV_X4 vscale_core_DW01_sub_6_U730 ( .A(pipeline_md_b[37]), .ZN(vscale_core_DW01_sub_6n425) );
  INV_X4 vscale_core_DW01_sub_6_U731 ( .A(pipeline_md_b[38]), .ZN(vscale_core_DW01_sub_6n424) );
  INV_X4 vscale_core_DW01_sub_6_U732 ( .A(pipeline_md_b[39]), .ZN(vscale_core_DW01_sub_6n423) );
  INV_X4 vscale_core_DW01_sub_6_U733 ( .A(pipeline_md_b[40]), .ZN(vscale_core_DW01_sub_6n422) );
  INV_X4 vscale_core_DW01_sub_6_U734 ( .A(pipeline_md_b[41]), .ZN(vscale_core_DW01_sub_6n421) );
  INV_X4 vscale_core_DW01_sub_6_U735 ( .A(pipeline_md_b[42]), .ZN(vscale_core_DW01_sub_6n420) );
  INV_X4 vscale_core_DW01_sub_6_U736 ( .A(pipeline_md_b[43]), .ZN(vscale_core_DW01_sub_6n419) );
  INV_X4 vscale_core_DW01_sub_6_U737 ( .A(pipeline_md_b[44]), .ZN(vscale_core_DW01_sub_6n418) );
  INV_X4 vscale_core_DW01_sub_6_U738 ( .A(pipeline_md_b[45]), .ZN(vscale_core_DW01_sub_6n417) );
  INV_X4 vscale_core_DW01_sub_6_U739 ( .A(pipeline_md_b[46]), .ZN(vscale_core_DW01_sub_6n416) );
  INV_X4 vscale_core_DW01_sub_6_U740 ( .A(pipeline_md_b[47]), .ZN(vscale_core_DW01_sub_6n415) );
  INV_X4 vscale_core_DW01_sub_6_U741 ( .A(pipeline_md_b[48]), .ZN(vscale_core_DW01_sub_6n414) );
  INV_X4 vscale_core_DW01_sub_6_U742 ( .A(pipeline_md_b[49]), .ZN(vscale_core_DW01_sub_6n413) );
  INV_X4 vscale_core_DW01_sub_6_U743 ( .A(pipeline_md_b[50]), .ZN(vscale_core_DW01_sub_6n412) );
  INV_X4 vscale_core_DW01_sub_6_U744 ( .A(pipeline_md_b[51]), .ZN(vscale_core_DW01_sub_6n411) );
  INV_X4 vscale_core_DW01_sub_6_U745 ( .A(pipeline_md_b[52]), .ZN(vscale_core_DW01_sub_6n410) );
  INV_X4 vscale_core_DW01_sub_6_U746 ( .A(pipeline_md_b[53]), .ZN(vscale_core_DW01_sub_6n409) );
  INV_X4 vscale_core_DW01_sub_6_U747 ( .A(pipeline_md_b[54]), .ZN(vscale_core_DW01_sub_6n408) );
  INV_X4 vscale_core_DW01_sub_6_U748 ( .A(pipeline_md_b[55]), .ZN(vscale_core_DW01_sub_6n407) );
  INV_X4 vscale_core_DW01_sub_6_U749 ( .A(pipeline_md_b[56]), .ZN(vscale_core_DW01_sub_6n406) );
  INV_X4 vscale_core_DW01_sub_6_U750 ( .A(pipeline_md_b[57]), .ZN(vscale_core_DW01_sub_6n405) );
  INV_X4 vscale_core_DW01_sub_6_U751 ( .A(pipeline_md_b[58]), .ZN(vscale_core_DW01_sub_6n404) );
  INV_X4 vscale_core_DW01_sub_6_U752 ( .A(pipeline_md_b[59]), .ZN(vscale_core_DW01_sub_6n403) );
  INV_X4 vscale_core_DW01_sub_6_U753 ( .A(pipeline_md_b[60]), .ZN(vscale_core_DW01_sub_6n402) );
  INV_X4 vscale_core_DW01_sub_6_U754 ( .A(pipeline_md_b[61]), .ZN(vscale_core_DW01_sub_6n401) );
  INV_X4 vscale_core_DW01_sub_6_U755 ( .A(pipeline_md_b[62]), .ZN(vscale_core_DW01_sub_6n400) );
  INV_X4 vscale_core_DW01_sub_6_U756 ( .A(vscale_core_DW01_sub_6n344), .ZN(vscale_core_DW01_sub_6n399) );
  INV_X4 vscale_core_DW01_sub_6_U757 ( .A(vscale_core_DW01_sub_6n340), .ZN(vscale_core_DW01_sub_6n398) );
  INV_X4 vscale_core_DW01_sub_6_U758 ( .A(vscale_core_DW01_sub_6n337), .ZN(vscale_core_DW01_sub_6n397) );
  INV_X4 vscale_core_DW01_sub_6_U759 ( .A(vscale_core_DW01_sub_6n326), .ZN(vscale_core_DW01_sub_6n395) );
  INV_X4 vscale_core_DW01_sub_6_U760 ( .A(vscale_core_DW01_sub_6n321), .ZN(vscale_core_DW01_sub_6n394) );
  INV_X4 vscale_core_DW01_sub_6_U761 ( .A(vscale_core_DW01_sub_6n318), .ZN(vscale_core_DW01_sub_6n393) );
  INV_X4 vscale_core_DW01_sub_6_U762 ( .A(vscale_core_DW01_sub_6n310), .ZN(vscale_core_DW01_sub_6n392) );
  INV_X4 vscale_core_DW01_sub_6_U763 ( .A(vscale_core_DW01_sub_6n307), .ZN(vscale_core_DW01_sub_6n391) );
  INV_X4 vscale_core_DW01_sub_6_U764 ( .A(vscale_core_DW01_sub_6n295), .ZN(vscale_core_DW01_sub_6n389) );
  INV_X4 vscale_core_DW01_sub_6_U765 ( .A(vscale_core_DW01_sub_6n282), .ZN(vscale_core_DW01_sub_6n387) );
  INV_X4 vscale_core_DW01_sub_6_U766 ( .A(vscale_core_DW01_sub_6n270), .ZN(vscale_core_DW01_sub_6n385) );
  INV_X4 vscale_core_DW01_sub_6_U767 ( .A(vscale_core_DW01_sub_6n255), .ZN(vscale_core_DW01_sub_6n383) );
  INV_X4 vscale_core_DW01_sub_6_U768 ( .A(vscale_core_DW01_sub_6n250), .ZN(vscale_core_DW01_sub_6n382) );
  INV_X4 vscale_core_DW01_sub_6_U769 ( .A(vscale_core_DW01_sub_6n247), .ZN(vscale_core_DW01_sub_6n381) );
  INV_X4 vscale_core_DW01_sub_6_U770 ( .A(vscale_core_DW01_sub_6n237), .ZN(vscale_core_DW01_sub_6n380) );
  INV_X4 vscale_core_DW01_sub_6_U771 ( .A(vscale_core_DW01_sub_6n234), .ZN(vscale_core_DW01_sub_6n379) );
  INV_X4 vscale_core_DW01_sub_6_U772 ( .A(vscale_core_DW01_sub_6n229), .ZN(vscale_core_DW01_sub_6n378) );
  INV_X4 vscale_core_DW01_sub_6_U773 ( .A(vscale_core_DW01_sub_6n226), .ZN(vscale_core_DW01_sub_6n377) );
  INV_X4 vscale_core_DW01_sub_6_U774 ( .A(vscale_core_DW01_sub_6n216), .ZN(vscale_core_DW01_sub_6n376) );
  INV_X4 vscale_core_DW01_sub_6_U775 ( .A(vscale_core_DW01_sub_6n213), .ZN(vscale_core_DW01_sub_6n375) );
  INV_X4 vscale_core_DW01_sub_6_U776 ( .A(vscale_core_DW01_sub_6n208), .ZN(vscale_core_DW01_sub_6n374) );
  INV_X4 vscale_core_DW01_sub_6_U777 ( .A(vscale_core_DW01_sub_6n205), .ZN(vscale_core_DW01_sub_6n373) );
  INV_X4 vscale_core_DW01_sub_6_U778 ( .A(vscale_core_DW01_sub_6n195), .ZN(vscale_core_DW01_sub_6n372) );
  INV_X4 vscale_core_DW01_sub_6_U779 ( .A(vscale_core_DW01_sub_6n192), .ZN(vscale_core_DW01_sub_6n371) );
  INV_X4 vscale_core_DW01_sub_6_U780 ( .A(vscale_core_DW01_sub_6n187), .ZN(vscale_core_DW01_sub_6n370) );
  INV_X4 vscale_core_DW01_sub_6_U781 ( .A(vscale_core_DW01_sub_6n184), .ZN(vscale_core_DW01_sub_6n369) );
  INV_X4 vscale_core_DW01_sub_6_U782 ( .A(vscale_core_DW01_sub_6n172), .ZN(vscale_core_DW01_sub_6n368) );
  INV_X4 vscale_core_DW01_sub_6_U783 ( .A(vscale_core_DW01_sub_6n169), .ZN(vscale_core_DW01_sub_6n367) );
  INV_X4 vscale_core_DW01_sub_6_U784 ( .A(vscale_core_DW01_sub_6n157), .ZN(vscale_core_DW01_sub_6n365) );
  INV_X4 vscale_core_DW01_sub_6_U785 ( .A(vscale_core_DW01_sub_6n144), .ZN(vscale_core_DW01_sub_6n363) );
  INV_X4 vscale_core_DW01_sub_6_U786 ( .A(vscale_core_DW01_sub_6n132), .ZN(vscale_core_DW01_sub_6n361) );
  INV_X4 vscale_core_DW01_sub_6_U787 ( .A(vscale_core_DW01_sub_6n116), .ZN(vscale_core_DW01_sub_6n359) );
  INV_X4 vscale_core_DW01_sub_6_U788 ( .A(vscale_core_DW01_sub_6n109), .ZN(vscale_core_DW01_sub_6n358) );
  INV_X4 vscale_core_DW01_sub_6_U789 ( .A(vscale_core_DW01_sub_6n104), .ZN(vscale_core_DW01_sub_6n357) );
  INV_X4 vscale_core_DW01_sub_6_U790 ( .A(vscale_core_DW01_sub_6n96), .ZN(vscale_core_DW01_sub_6n355) );
  INV_X4 vscale_core_DW01_sub_6_U791 ( .A(vscale_core_DW01_sub_6n88), .ZN(vscale_core_DW01_sub_6n353) );
  INV_X4 vscale_core_DW01_sub_6_U792 ( .A(vscale_core_DW01_sub_6n80), .ZN(vscale_core_DW01_sub_6n351) );
  INV_X4 vscale_core_DW01_sub_6_U793 ( .A(vscale_core_DW01_sub_6n72), .ZN(vscale_core_DW01_sub_6n349) );
  INV_X4 vscale_core_DW01_sub_6_U794 ( .A(vscale_core_DW01_sub_6n64), .ZN(vscale_core_DW01_sub_6n347) );
  INV_X4 vscale_core_DW01_sub_6_U795 ( .A(vscale_core_DW01_sub_6n343), .ZN(vscale_core_DW01_sub_6n342) );
  INV_X4 vscale_core_DW01_sub_6_U796 ( .A(vscale_core_DW01_sub_6n334), .ZN(vscale_core_DW01_sub_6n333) );
  INV_X4 vscale_core_DW01_sub_6_U797 ( .A(vscale_core_DW01_sub_6n332), .ZN(vscale_core_DW01_sub_6n330) );
  INV_X4 vscale_core_DW01_sub_6_U798 ( .A(vscale_core_DW01_sub_6n331), .ZN(vscale_core_DW01_sub_6n396) );
  INV_X4 vscale_core_DW01_sub_6_U799 ( .A(vscale_core_DW01_sub_6n313), .ZN(vscale_core_DW01_sub_6n312) );
  INV_X4 vscale_core_DW01_sub_6_U800 ( .A(vscale_core_DW01_sub_6n306), .ZN(vscale_core_DW01_sub_6n304) );
  INV_X4 vscale_core_DW01_sub_6_U801 ( .A(vscale_core_DW01_sub_6n305), .ZN(vscale_core_DW01_sub_6n303) );
  INV_X4 vscale_core_DW01_sub_6_U802 ( .A(vscale_core_DW01_sub_6n301), .ZN(vscale_core_DW01_sub_6n299) );
  INV_X4 vscale_core_DW01_sub_6_U803 ( .A(vscale_core_DW01_sub_6n300), .ZN(vscale_core_DW01_sub_6n390) );
  INV_X4 vscale_core_DW01_sub_6_U804 ( .A(vscale_core_DW01_sub_6n290), .ZN(vscale_core_DW01_sub_6n289) );
  INV_X4 vscale_core_DW01_sub_6_U805 ( .A(vscale_core_DW01_sub_6n288), .ZN(vscale_core_DW01_sub_6n286) );
  INV_X4 vscale_core_DW01_sub_6_U806 ( .A(vscale_core_DW01_sub_6n287), .ZN(vscale_core_DW01_sub_6n388) );
  INV_X4 vscale_core_DW01_sub_6_U807 ( .A(vscale_core_DW01_sub_6n281), .ZN(vscale_core_DW01_sub_6n279) );
  INV_X4 vscale_core_DW01_sub_6_U808 ( .A(vscale_core_DW01_sub_6n280), .ZN(vscale_core_DW01_sub_6n278) );
  INV_X4 vscale_core_DW01_sub_6_U809 ( .A(vscale_core_DW01_sub_6n276), .ZN(vscale_core_DW01_sub_6n274) );
  INV_X4 vscale_core_DW01_sub_6_U810 ( .A(vscale_core_DW01_sub_6n275), .ZN(vscale_core_DW01_sub_6n386) );
  INV_X4 vscale_core_DW01_sub_6_U811 ( .A(vscale_core_DW01_sub_6n263), .ZN(vscale_core_DW01_sub_6n262) );
  INV_X4 vscale_core_DW01_sub_6_U812 ( .A(vscale_core_DW01_sub_6n261), .ZN(vscale_core_DW01_sub_6n259) );
  INV_X4 vscale_core_DW01_sub_6_U813 ( .A(vscale_core_DW01_sub_6n260), .ZN(vscale_core_DW01_sub_6n384) );
  INV_X4 vscale_core_DW01_sub_6_U814 ( .A(vscale_core_DW01_sub_6n244), .ZN(vscale_core_DW01_sub_6n242) );
  INV_X4 vscale_core_DW01_sub_6_U815 ( .A(vscale_core_DW01_sub_6n243), .ZN(vscale_core_DW01_sub_6n241) );
  INV_X4 vscale_core_DW01_sub_6_U816 ( .A(vscale_core_DW01_sub_6n240), .ZN(vscale_core_DW01_sub_6n239) );
  INV_X4 vscale_core_DW01_sub_6_U817 ( .A(vscale_core_DW01_sub_6n219), .ZN(vscale_core_DW01_sub_6n218) );
  INV_X4 vscale_core_DW01_sub_6_U818 ( .A(vscale_core_DW01_sub_6n202), .ZN(vscale_core_DW01_sub_6n200) );
  INV_X4 vscale_core_DW01_sub_6_U819 ( .A(vscale_core_DW01_sub_6n201), .ZN(vscale_core_DW01_sub_6n199) );
  INV_X4 vscale_core_DW01_sub_6_U820 ( .A(vscale_core_DW01_sub_6n198), .ZN(vscale_core_DW01_sub_6n197) );
  INV_X4 vscale_core_DW01_sub_6_U821 ( .A(vscale_core_DW01_sub_6n175), .ZN(vscale_core_DW01_sub_6n174) );
  INV_X4 vscale_core_DW01_sub_6_U822 ( .A(vscale_core_DW01_sub_6n168), .ZN(vscale_core_DW01_sub_6n166) );
  INV_X4 vscale_core_DW01_sub_6_U823 ( .A(vscale_core_DW01_sub_6n167), .ZN(vscale_core_DW01_sub_6n165) );
  INV_X4 vscale_core_DW01_sub_6_U824 ( .A(vscale_core_DW01_sub_6n163), .ZN(vscale_core_DW01_sub_6n161) );
  INV_X4 vscale_core_DW01_sub_6_U825 ( .A(vscale_core_DW01_sub_6n162), .ZN(vscale_core_DW01_sub_6n366) );
  INV_X4 vscale_core_DW01_sub_6_U826 ( .A(vscale_core_DW01_sub_6n152), .ZN(vscale_core_DW01_sub_6n151) );
  INV_X4 vscale_core_DW01_sub_6_U827 ( .A(vscale_core_DW01_sub_6n150), .ZN(vscale_core_DW01_sub_6n148) );
  INV_X4 vscale_core_DW01_sub_6_U828 ( .A(vscale_core_DW01_sub_6n149), .ZN(vscale_core_DW01_sub_6n364) );
  INV_X4 vscale_core_DW01_sub_6_U829 ( .A(vscale_core_DW01_sub_6n143), .ZN(vscale_core_DW01_sub_6n141) );
  INV_X4 vscale_core_DW01_sub_6_U830 ( .A(vscale_core_DW01_sub_6n142), .ZN(vscale_core_DW01_sub_6n140) );
  INV_X4 vscale_core_DW01_sub_6_U831 ( .A(vscale_core_DW01_sub_6n138), .ZN(vscale_core_DW01_sub_6n136) );
  INV_X4 vscale_core_DW01_sub_6_U832 ( .A(vscale_core_DW01_sub_6n137), .ZN(vscale_core_DW01_sub_6n362) );
  INV_X4 vscale_core_DW01_sub_6_U833 ( .A(vscale_core_DW01_sub_6n127), .ZN(vscale_core_DW01_sub_6n125) );
  INV_X4 vscale_core_DW01_sub_6_U834 ( .A(vscale_core_DW01_sub_6n126), .ZN(vscale_core_DW01_sub_6n124) );
  INV_X4 vscale_core_DW01_sub_6_U835 ( .A(vscale_core_DW01_sub_6n122), .ZN(vscale_core_DW01_sub_6n120) );
  INV_X4 vscale_core_DW01_sub_6_U836 ( .A(vscale_core_DW01_sub_6n121), .ZN(vscale_core_DW01_sub_6n360) );
  INV_X4 vscale_core_DW01_sub_6_U837 ( .A(vscale_core_DW01_sub_6n102), .ZN(vscale_core_DW01_sub_6n100) );
;
  vscale_core_DW01_add_5 pipeline_md_add_104 

  XOR2_X2 vscale_core_DW01_add_5_U1 ( .A(n10234), .B(vscale_core_DW01_add_5n55), .Z(pipeline_md_N249) );
  FA_X1 vscale_core_DW01_add_5_U2 ( .A(pipeline_md_b[62]), .B(pipeline_md_result[62]), .CI(vscale_core_DW01_add_5n56), .CO(vscale_core_DW01_add_5n55), .S(pipeline_md_N248) );
  FA_X1 vscale_core_DW01_add_5_U3 ( .A(pipeline_md_b[61]), .B(pipeline_md_result[61]), .CI(vscale_core_DW01_add_5n57), .CO(vscale_core_DW01_add_5n56), .S(pipeline_md_N247) );
  FA_X1 vscale_core_DW01_add_5_U4 ( .A(pipeline_md_b[60]), .B(pipeline_md_result[60]), .CI(vscale_core_DW01_add_5n58), .CO(vscale_core_DW01_add_5n57), .S(pipeline_md_N246) );
  FA_X1 vscale_core_DW01_add_5_U5 ( .A(pipeline_md_b[59]), .B(pipeline_md_result[59]), .CI(vscale_core_DW01_add_5n59), .CO(vscale_core_DW01_add_5n58), .S(pipeline_md_N245) );
  FA_X1 vscale_core_DW01_add_5_U6 ( .A(pipeline_md_b[58]), .B(pipeline_md_result[58]), .CI(vscale_core_DW01_add_5n60), .CO(vscale_core_DW01_add_5n59), .S(pipeline_md_N244) );
  FA_X1 vscale_core_DW01_add_5_U7 ( .A(pipeline_md_b[57]), .B(pipeline_md_result[57]), .CI(vscale_core_DW01_add_5n61), .CO(vscale_core_DW01_add_5n60), .S(pipeline_md_N243) );
  FA_X1 vscale_core_DW01_add_5_U8 ( .A(pipeline_md_b[56]), .B(pipeline_md_result[56]), .CI(vscale_core_DW01_add_5n62), .CO(vscale_core_DW01_add_5n61), .S(pipeline_md_N242) );
  FA_X1 vscale_core_DW01_add_5_U9 ( .A(pipeline_md_b[55]), .B(pipeline_md_result[55]), .CI(vscale_core_DW01_add_5n63), .CO(vscale_core_DW01_add_5n62), .S(pipeline_md_N241) );
  FA_X1 vscale_core_DW01_add_5_U10 ( .A(pipeline_md_b[54]), .B(pipeline_md_result[54]), .CI(vscale_core_DW01_add_5n64), .CO(vscale_core_DW01_add_5n63), .S(pipeline_md_N240) );
  XOR2_X2 vscale_core_DW01_add_5_U11 ( .A(vscale_core_DW01_add_5n1), .B(vscale_core_DW01_add_5n67), .Z(pipeline_md_N239) );
  NAND2_X2 vscale_core_DW01_add_5_U13 ( .A1(vscale_core_DW01_add_5n349), .A2(vscale_core_DW01_add_5n66), .ZN(vscale_core_DW01_add_5n1) );
  NAND2_X2 vscale_core_DW01_add_5_U16 ( .A1(pipeline_md_b[53]), .A2(pipeline_md_result[53]), .ZN(vscale_core_DW01_add_5n66) );
  XNOR2_X2 vscale_core_DW01_add_5_U17 ( .A(vscale_core_DW01_add_5n72), .B(vscale_core_DW01_add_5n2), .ZN(pipeline_md_N238) );
  NAND2_X2 vscale_core_DW01_add_5_U21 ( .A1(vscale_core_DW01_add_5n606), .A2(vscale_core_DW01_add_5n71), .ZN(vscale_core_DW01_add_5n2) );
  NAND2_X2 vscale_core_DW01_add_5_U24 ( .A1(pipeline_md_b[52]), .A2(pipeline_md_result[52]), .ZN(vscale_core_DW01_add_5n71) );
  XOR2_X2 vscale_core_DW01_add_5_U25 ( .A(vscale_core_DW01_add_5n3), .B(vscale_core_DW01_add_5n75), .Z(pipeline_md_N237) );
  NAND2_X2 vscale_core_DW01_add_5_U27 ( .A1(vscale_core_DW01_add_5n351), .A2(vscale_core_DW01_add_5n74), .ZN(vscale_core_DW01_add_5n3) );
  NAND2_X2 vscale_core_DW01_add_5_U30 ( .A1(pipeline_md_b[51]), .A2(pipeline_md_result[51]), .ZN(vscale_core_DW01_add_5n74) );
  XNOR2_X2 vscale_core_DW01_add_5_U31 ( .A(vscale_core_DW01_add_5n80), .B(vscale_core_DW01_add_5n4), .ZN(pipeline_md_N236) );
  NAND2_X2 vscale_core_DW01_add_5_U35 ( .A1(vscale_core_DW01_add_5n603), .A2(vscale_core_DW01_add_5n79), .ZN(vscale_core_DW01_add_5n4) );
  NAND2_X2 vscale_core_DW01_add_5_U38 ( .A1(pipeline_md_b[50]), .A2(pipeline_md_result[50]), .ZN(vscale_core_DW01_add_5n79) );
  XOR2_X2 vscale_core_DW01_add_5_U39 ( .A(vscale_core_DW01_add_5n5), .B(vscale_core_DW01_add_5n83), .Z(pipeline_md_N235) );
  NAND2_X2 vscale_core_DW01_add_5_U41 ( .A1(vscale_core_DW01_add_5n353), .A2(vscale_core_DW01_add_5n82), .ZN(vscale_core_DW01_add_5n5) );
  NAND2_X2 vscale_core_DW01_add_5_U44 ( .A1(pipeline_md_b[49]), .A2(pipeline_md_result[49]), .ZN(vscale_core_DW01_add_5n82) );
  XNOR2_X2 vscale_core_DW01_add_5_U45 ( .A(vscale_core_DW01_add_5n88), .B(vscale_core_DW01_add_5n6), .ZN(pipeline_md_N234) );
  NAND2_X2 vscale_core_DW01_add_5_U49 ( .A1(vscale_core_DW01_add_5n605), .A2(vscale_core_DW01_add_5n87), .ZN(vscale_core_DW01_add_5n6) );
  NAND2_X2 vscale_core_DW01_add_5_U52 ( .A1(pipeline_md_b[48]), .A2(pipeline_md_result[48]), .ZN(vscale_core_DW01_add_5n87) );
  XOR2_X2 vscale_core_DW01_add_5_U53 ( .A(vscale_core_DW01_add_5n7), .B(vscale_core_DW01_add_5n91), .Z(pipeline_md_N233) );
  NAND2_X2 vscale_core_DW01_add_5_U55 ( .A1(vscale_core_DW01_add_5n355), .A2(vscale_core_DW01_add_5n90), .ZN(vscale_core_DW01_add_5n7) );
  NAND2_X2 vscale_core_DW01_add_5_U58 ( .A1(pipeline_md_b[47]), .A2(pipeline_md_result[47]), .ZN(vscale_core_DW01_add_5n90) );
  XNOR2_X2 vscale_core_DW01_add_5_U59 ( .A(vscale_core_DW01_add_5n96), .B(vscale_core_DW01_add_5n8), .ZN(pipeline_md_N232) );
  NAND2_X2 vscale_core_DW01_add_5_U63 ( .A1(vscale_core_DW01_add_5n604), .A2(vscale_core_DW01_add_5n95), .ZN(vscale_core_DW01_add_5n8) );
  NAND2_X2 vscale_core_DW01_add_5_U66 ( .A1(pipeline_md_b[46]), .A2(pipeline_md_result[46]), .ZN(vscale_core_DW01_add_5n95) );
  XOR2_X2 vscale_core_DW01_add_5_U67 ( .A(vscale_core_DW01_add_5n9), .B(vscale_core_DW01_add_5n99), .Z(pipeline_md_N231) );
  NAND2_X2 vscale_core_DW01_add_5_U69 ( .A1(vscale_core_DW01_add_5n357), .A2(vscale_core_DW01_add_5n98), .ZN(vscale_core_DW01_add_5n9) );
  NAND2_X2 vscale_core_DW01_add_5_U72 ( .A1(pipeline_md_b[45]), .A2(pipeline_md_result[45]), .ZN(vscale_core_DW01_add_5n98) );
  XNOR2_X2 vscale_core_DW01_add_5_U73 ( .A(vscale_core_DW01_add_5n104), .B(vscale_core_DW01_add_5n10), .ZN(pipeline_md_N230) );
  NAND2_X2 vscale_core_DW01_add_5_U77 ( .A1(vscale_core_DW01_add_5n602), .A2(vscale_core_DW01_add_5n103), .ZN(vscale_core_DW01_add_5n10) );
  NAND2_X2 vscale_core_DW01_add_5_U80 ( .A1(pipeline_md_b[44]), .A2(pipeline_md_result[44]), .ZN(vscale_core_DW01_add_5n103) );
  XOR2_X2 vscale_core_DW01_add_5_U81 ( .A(vscale_core_DW01_add_5n11), .B(vscale_core_DW01_add_5n107), .Z(pipeline_md_N229) );
  NAND2_X2 vscale_core_DW01_add_5_U83 ( .A1(vscale_core_DW01_add_5n359), .A2(vscale_core_DW01_add_5n106), .ZN(vscale_core_DW01_add_5n11) );
  NAND2_X2 vscale_core_DW01_add_5_U86 ( .A1(pipeline_md_b[43]), .A2(pipeline_md_result[43]), .ZN(vscale_core_DW01_add_5n106) );
  XNOR2_X2 vscale_core_DW01_add_5_U87 ( .A(vscale_core_DW01_add_5n112), .B(vscale_core_DW01_add_5n12), .ZN(pipeline_md_N228) );
  NAND2_X2 vscale_core_DW01_add_5_U91 ( .A1(vscale_core_DW01_add_5n360), .A2(vscale_core_DW01_add_5n111), .ZN(vscale_core_DW01_add_5n12) );
  NAND2_X2 vscale_core_DW01_add_5_U94 ( .A1(pipeline_md_b[42]), .A2(pipeline_md_result[42]), .ZN(vscale_core_DW01_add_5n111) );
  XOR2_X2 vscale_core_DW01_add_5_U95 ( .A(vscale_core_DW01_add_5n13), .B(vscale_core_DW01_add_5n119), .Z(pipeline_md_N227) );
  NAND2_X2 vscale_core_DW01_add_5_U97 ( .A1(vscale_core_DW01_add_5n127), .A2(vscale_core_DW01_add_5n115), .ZN(vscale_core_DW01_add_5n113) );
  NAND2_X2 vscale_core_DW01_add_5_U101 ( .A1(vscale_core_DW01_add_5n361), .A2(vscale_core_DW01_add_5n118), .ZN(vscale_core_DW01_add_5n13) );
  NAND2_X2 vscale_core_DW01_add_5_U104 ( .A1(pipeline_md_b[41]), .A2(pipeline_md_result[41]), .ZN(vscale_core_DW01_add_5n118) );
  XNOR2_X2 vscale_core_DW01_add_5_U105 ( .A(vscale_core_DW01_add_5n124), .B(vscale_core_DW01_add_5n14), .ZN(pipeline_md_N226) );
  NAND2_X2 vscale_core_DW01_add_5_U109 ( .A1(vscale_core_DW01_add_5n362), .A2(vscale_core_DW01_add_5n123), .ZN(vscale_core_DW01_add_5n14) );
  NAND2_X2 vscale_core_DW01_add_5_U112 ( .A1(pipeline_md_b[40]), .A2(pipeline_md_result[40]), .ZN(vscale_core_DW01_add_5n123) );
  XOR2_X2 vscale_core_DW01_add_5_U113 ( .A(vscale_core_DW01_add_5n15), .B(vscale_core_DW01_add_5n135), .Z(pipeline_md_N225) );
  NAND2_X2 vscale_core_DW01_add_5_U119 ( .A1(vscale_core_DW01_add_5n143), .A2(vscale_core_DW01_add_5n131), .ZN(vscale_core_DW01_add_5n129) );
  NAND2_X2 vscale_core_DW01_add_5_U123 ( .A1(vscale_core_DW01_add_5n363), .A2(vscale_core_DW01_add_5n134), .ZN(vscale_core_DW01_add_5n15) );
  NAND2_X2 vscale_core_DW01_add_5_U126 ( .A1(pipeline_md_b[39]), .A2(pipeline_md_result[39]), .ZN(vscale_core_DW01_add_5n134) );
  XNOR2_X2 vscale_core_DW01_add_5_U127 ( .A(vscale_core_DW01_add_5n140), .B(vscale_core_DW01_add_5n16), .ZN(pipeline_md_N224) );
  NAND2_X2 vscale_core_DW01_add_5_U131 ( .A1(vscale_core_DW01_add_5n364), .A2(vscale_core_DW01_add_5n139), .ZN(vscale_core_DW01_add_5n16) );
  NAND2_X2 vscale_core_DW01_add_5_U134 ( .A1(pipeline_md_b[38]), .A2(pipeline_md_result[38]), .ZN(vscale_core_DW01_add_5n139) );
  XOR2_X2 vscale_core_DW01_add_5_U135 ( .A(vscale_core_DW01_add_5n17), .B(vscale_core_DW01_add_5n147), .Z(pipeline_md_N223) );
  NAND2_X2 vscale_core_DW01_add_5_U141 ( .A1(vscale_core_DW01_add_5n365), .A2(vscale_core_DW01_add_5n146), .ZN(vscale_core_DW01_add_5n17) );
  NAND2_X2 vscale_core_DW01_add_5_U144 ( .A1(pipeline_md_b[37]), .A2(pipeline_md_result[37]), .ZN(vscale_core_DW01_add_5n146) );
  XOR2_X2 vscale_core_DW01_add_5_U145 ( .A(vscale_core_DW01_add_5n18), .B(vscale_core_DW01_add_5n152), .Z(pipeline_md_N222) );
  NAND2_X2 vscale_core_DW01_add_5_U149 ( .A1(vscale_core_DW01_add_5n366), .A2(vscale_core_DW01_add_5n151), .ZN(vscale_core_DW01_add_5n18) );
  NAND2_X2 vscale_core_DW01_add_5_U152 ( .A1(pipeline_md_b[36]), .A2(pipeline_md_result[36]), .ZN(vscale_core_DW01_add_5n151) );
  XOR2_X2 vscale_core_DW01_add_5_U153 ( .A(vscale_core_DW01_add_5n19), .B(vscale_core_DW01_add_5n160), .Z(pipeline_md_N221) );
  NAND2_X2 vscale_core_DW01_add_5_U156 ( .A1(vscale_core_DW01_add_5n168), .A2(vscale_core_DW01_add_5n156), .ZN(vscale_core_DW01_add_5n154) );
  NAND2_X2 vscale_core_DW01_add_5_U160 ( .A1(vscale_core_DW01_add_5n367), .A2(vscale_core_DW01_add_5n159), .ZN(vscale_core_DW01_add_5n19) );
  NAND2_X2 vscale_core_DW01_add_5_U163 ( .A1(pipeline_md_b[35]), .A2(pipeline_md_result[35]), .ZN(vscale_core_DW01_add_5n159) );
  XNOR2_X2 vscale_core_DW01_add_5_U164 ( .A(vscale_core_DW01_add_5n165), .B(vscale_core_DW01_add_5n20), .ZN(pipeline_md_N220) );
  NAND2_X2 vscale_core_DW01_add_5_U168 ( .A1(vscale_core_DW01_add_5n368), .A2(vscale_core_DW01_add_5n164), .ZN(vscale_core_DW01_add_5n20) );
  NAND2_X2 vscale_core_DW01_add_5_U171 ( .A1(pipeline_md_b[34]), .A2(pipeline_md_result[34]), .ZN(vscale_core_DW01_add_5n164) );
  XNOR2_X2 vscale_core_DW01_add_5_U172 ( .A(vscale_core_DW01_add_5n172), .B(vscale_core_DW01_add_5n21), .ZN(pipeline_md_N219) );
  NAND2_X2 vscale_core_DW01_add_5_U178 ( .A1(vscale_core_DW01_add_5n369), .A2(vscale_core_DW01_add_5n171), .ZN(vscale_core_DW01_add_5n21) );
  NAND2_X2 vscale_core_DW01_add_5_U181 ( .A1(pipeline_md_b[33]), .A2(pipeline_md_result[33]), .ZN(vscale_core_DW01_add_5n171) );
  XOR2_X2 vscale_core_DW01_add_5_U182 ( .A(vscale_core_DW01_add_5n22), .B(vscale_core_DW01_add_5n175), .Z(pipeline_md_N218) );
  NAND2_X2 vscale_core_DW01_add_5_U184 ( .A1(vscale_core_DW01_add_5n370), .A2(vscale_core_DW01_add_5n174), .ZN(vscale_core_DW01_add_5n22) );
  NAND2_X2 vscale_core_DW01_add_5_U187 ( .A1(pipeline_md_b[32]), .A2(pipeline_md_result[32]), .ZN(vscale_core_DW01_add_5n174) );
  XNOR2_X2 vscale_core_DW01_add_5_U188 ( .A(vscale_core_DW01_add_5n187), .B(vscale_core_DW01_add_5n23), .ZN(pipeline_md_N217) );
  NAND2_X2 vscale_core_DW01_add_5_U191 ( .A1(vscale_core_DW01_add_5n221), .A2(vscale_core_DW01_add_5n179), .ZN(vscale_core_DW01_add_5n177) );
  NAND2_X2 vscale_core_DW01_add_5_U195 ( .A1(vscale_core_DW01_add_5n191), .A2(vscale_core_DW01_add_5n183), .ZN(vscale_core_DW01_add_5n181) );
  NAND2_X2 vscale_core_DW01_add_5_U199 ( .A1(vscale_core_DW01_add_5n371), .A2(vscale_core_DW01_add_5n186), .ZN(vscale_core_DW01_add_5n23) );
  NAND2_X2 vscale_core_DW01_add_5_U202 ( .A1(pipeline_md_b[31]), .A2(pipeline_md_resp_result[31]), .ZN(vscale_core_DW01_add_5n186) );
  XOR2_X2 vscale_core_DW01_add_5_U203 ( .A(vscale_core_DW01_add_5n24), .B(vscale_core_DW01_add_5n190), .Z(pipeline_md_N216) );
  NAND2_X2 vscale_core_DW01_add_5_U205 ( .A1(vscale_core_DW01_add_5n372), .A2(vscale_core_DW01_add_5n189), .ZN(vscale_core_DW01_add_5n24) );
  NAND2_X2 vscale_core_DW01_add_5_U208 ( .A1(pipeline_md_b[30]), .A2(pipeline_md_resp_result[30]), .ZN(vscale_core_DW01_add_5n189) );
  XNOR2_X2 vscale_core_DW01_add_5_U209 ( .A(vscale_core_DW01_add_5n195), .B(vscale_core_DW01_add_5n25), .ZN(pipeline_md_N215) );
  NAND2_X2 vscale_core_DW01_add_5_U213 ( .A1(vscale_core_DW01_add_5n373), .A2(vscale_core_DW01_add_5n194), .ZN(vscale_core_DW01_add_5n25) );
  NAND2_X2 vscale_core_DW01_add_5_U216 ( .A1(pipeline_md_b[29]), .A2(pipeline_md_resp_result[29]), .ZN(vscale_core_DW01_add_5n194) );
  XNOR2_X2 vscale_core_DW01_add_5_U217 ( .A(vscale_core_DW01_add_5n198), .B(vscale_core_DW01_add_5n26), .ZN(pipeline_md_N214) );
  NAND2_X2 vscale_core_DW01_add_5_U219 ( .A1(vscale_core_DW01_add_5n374), .A2(vscale_core_DW01_add_5n197), .ZN(vscale_core_DW01_add_5n26) );
  NAND2_X2 vscale_core_DW01_add_5_U222 ( .A1(pipeline_md_b[28]), .A2(pipeline_md_resp_result[28]), .ZN(vscale_core_DW01_add_5n197) );
  XNOR2_X2 vscale_core_DW01_add_5_U223 ( .A(vscale_core_DW01_add_5n208), .B(vscale_core_DW01_add_5n27), .ZN(pipeline_md_N213) );
  NAND2_X2 vscale_core_DW01_add_5_U228 ( .A1(vscale_core_DW01_add_5n212), .A2(vscale_core_DW01_add_5n204), .ZN(vscale_core_DW01_add_5n202) );
  NAND2_X2 vscale_core_DW01_add_5_U232 ( .A1(vscale_core_DW01_add_5n375), .A2(vscale_core_DW01_add_5n207), .ZN(vscale_core_DW01_add_5n27) );
  NAND2_X2 vscale_core_DW01_add_5_U235 ( .A1(pipeline_md_b[27]), .A2(pipeline_md_resp_result[27]), .ZN(vscale_core_DW01_add_5n207) );
  XOR2_X2 vscale_core_DW01_add_5_U236 ( .A(vscale_core_DW01_add_5n28), .B(vscale_core_DW01_add_5n211), .Z(pipeline_md_N212) );
  NAND2_X2 vscale_core_DW01_add_5_U238 ( .A1(vscale_core_DW01_add_5n376), .A2(vscale_core_DW01_add_5n210), .ZN(vscale_core_DW01_add_5n28) );
  NAND2_X2 vscale_core_DW01_add_5_U241 ( .A1(pipeline_md_b[26]), .A2(pipeline_md_resp_result[26]), .ZN(vscale_core_DW01_add_5n210) );
  XNOR2_X2 vscale_core_DW01_add_5_U242 ( .A(vscale_core_DW01_add_5n216), .B(vscale_core_DW01_add_5n29), .ZN(pipeline_md_N211) );
  NAND2_X2 vscale_core_DW01_add_5_U246 ( .A1(vscale_core_DW01_add_5n377), .A2(vscale_core_DW01_add_5n215), .ZN(vscale_core_DW01_add_5n29) );
  NAND2_X2 vscale_core_DW01_add_5_U249 ( .A1(pipeline_md_b[25]), .A2(pipeline_md_resp_result[25]), .ZN(vscale_core_DW01_add_5n215) );
  XNOR2_X2 vscale_core_DW01_add_5_U250 ( .A(vscale_core_DW01_add_5n219), .B(vscale_core_DW01_add_5n30), .ZN(pipeline_md_N210) );
  NAND2_X2 vscale_core_DW01_add_5_U252 ( .A1(vscale_core_DW01_add_5n378), .A2(vscale_core_DW01_add_5n218), .ZN(vscale_core_DW01_add_5n30) );
  NAND2_X2 vscale_core_DW01_add_5_U255 ( .A1(pipeline_md_b[24]), .A2(pipeline_md_resp_result[24]), .ZN(vscale_core_DW01_add_5n218) );
  XNOR2_X2 vscale_core_DW01_add_5_U256 ( .A(vscale_core_DW01_add_5n229), .B(vscale_core_DW01_add_5n31), .ZN(pipeline_md_N209) );
  NAND2_X2 vscale_core_DW01_add_5_U261 ( .A1(vscale_core_DW01_add_5n233), .A2(vscale_core_DW01_add_5n225), .ZN(vscale_core_DW01_add_5n223) );
  NAND2_X2 vscale_core_DW01_add_5_U265 ( .A1(vscale_core_DW01_add_5n379), .A2(vscale_core_DW01_add_5n228), .ZN(vscale_core_DW01_add_5n31) );
  NAND2_X2 vscale_core_DW01_add_5_U268 ( .A1(pipeline_md_b[23]), .A2(pipeline_md_resp_result[23]), .ZN(vscale_core_DW01_add_5n228) );
  XOR2_X2 vscale_core_DW01_add_5_U269 ( .A(vscale_core_DW01_add_5n32), .B(vscale_core_DW01_add_5n232), .Z(pipeline_md_N208) );
  NAND2_X2 vscale_core_DW01_add_5_U271 ( .A1(vscale_core_DW01_add_5n380), .A2(vscale_core_DW01_add_5n231), .ZN(vscale_core_DW01_add_5n32) );
  NAND2_X2 vscale_core_DW01_add_5_U274 ( .A1(pipeline_md_b[22]), .A2(pipeline_md_resp_result[22]), .ZN(vscale_core_DW01_add_5n231) );
  XNOR2_X2 vscale_core_DW01_add_5_U275 ( .A(vscale_core_DW01_add_5n237), .B(vscale_core_DW01_add_5n33), .ZN(pipeline_md_N207) );
  NAND2_X2 vscale_core_DW01_add_5_U279 ( .A1(vscale_core_DW01_add_5n381), .A2(vscale_core_DW01_add_5n236), .ZN(vscale_core_DW01_add_5n33) );
  NAND2_X2 vscale_core_DW01_add_5_U282 ( .A1(pipeline_md_b[21]), .A2(pipeline_md_resp_result[21]), .ZN(vscale_core_DW01_add_5n236) );
  XNOR2_X2 vscale_core_DW01_add_5_U283 ( .A(vscale_core_DW01_add_5n240), .B(vscale_core_DW01_add_5n34), .ZN(pipeline_md_N206) );
  NAND2_X2 vscale_core_DW01_add_5_U285 ( .A1(vscale_core_DW01_add_5n382), .A2(vscale_core_DW01_add_5n239), .ZN(vscale_core_DW01_add_5n34) );
  NAND2_X2 vscale_core_DW01_add_5_U288 ( .A1(pipeline_md_b[20]), .A2(pipeline_md_resp_result[20]), .ZN(vscale_core_DW01_add_5n239) );
  XNOR2_X2 vscale_core_DW01_add_5_U289 ( .A(vscale_core_DW01_add_5n250), .B(vscale_core_DW01_add_5n35), .ZN(pipeline_md_N205) );
  NAND2_X2 vscale_core_DW01_add_5_U294 ( .A1(vscale_core_DW01_add_5n254), .A2(vscale_core_DW01_add_5n246), .ZN(vscale_core_DW01_add_5n244) );
  NAND2_X2 vscale_core_DW01_add_5_U298 ( .A1(vscale_core_DW01_add_5n383), .A2(vscale_core_DW01_add_5n249), .ZN(vscale_core_DW01_add_5n35) );
  NAND2_X2 vscale_core_DW01_add_5_U301 ( .A1(pipeline_md_b[19]), .A2(pipeline_md_resp_result[19]), .ZN(vscale_core_DW01_add_5n249) );
  XOR2_X2 vscale_core_DW01_add_5_U302 ( .A(vscale_core_DW01_add_5n36), .B(vscale_core_DW01_add_5n253), .Z(pipeline_md_N204) );
  NAND2_X2 vscale_core_DW01_add_5_U304 ( .A1(vscale_core_DW01_add_5n384), .A2(vscale_core_DW01_add_5n252), .ZN(vscale_core_DW01_add_5n36) );
  NAND2_X2 vscale_core_DW01_add_5_U307 ( .A1(pipeline_md_b[18]), .A2(pipeline_md_resp_result[18]), .ZN(vscale_core_DW01_add_5n252) );
  XOR2_X2 vscale_core_DW01_add_5_U308 ( .A(vscale_core_DW01_add_5n37), .B(vscale_core_DW01_add_5n258), .Z(pipeline_md_N203) );
  NAND2_X2 vscale_core_DW01_add_5_U312 ( .A1(vscale_core_DW01_add_5n385), .A2(vscale_core_DW01_add_5n257), .ZN(vscale_core_DW01_add_5n37) );
  NAND2_X2 vscale_core_DW01_add_5_U315 ( .A1(pipeline_md_b[17]), .A2(pipeline_md_resp_result[17]), .ZN(vscale_core_DW01_add_5n257) );
  XNOR2_X2 vscale_core_DW01_add_5_U316 ( .A(vscale_core_DW01_add_5n263), .B(vscale_core_DW01_add_5n38), .ZN(pipeline_md_N202) );
  NAND2_X2 vscale_core_DW01_add_5_U320 ( .A1(vscale_core_DW01_add_5n386), .A2(vscale_core_DW01_add_5n262), .ZN(vscale_core_DW01_add_5n38) );
  NAND2_X2 vscale_core_DW01_add_5_U323 ( .A1(pipeline_md_b[16]), .A2(pipeline_md_resp_result[16]), .ZN(vscale_core_DW01_add_5n262) );
  XOR2_X2 vscale_core_DW01_add_5_U324 ( .A(vscale_core_DW01_add_5n39), .B(vscale_core_DW01_add_5n273), .Z(pipeline_md_N201) );
  NAND2_X2 vscale_core_DW01_add_5_U329 ( .A1(vscale_core_DW01_add_5n281), .A2(vscale_core_DW01_add_5n269), .ZN(vscale_core_DW01_add_5n267) );
  NAND2_X2 vscale_core_DW01_add_5_U333 ( .A1(vscale_core_DW01_add_5n387), .A2(vscale_core_DW01_add_5n272), .ZN(vscale_core_DW01_add_5n39) );
  NAND2_X2 vscale_core_DW01_add_5_U336 ( .A1(pipeline_md_b[15]), .A2(pipeline_md_resp_result[15]), .ZN(vscale_core_DW01_add_5n272) );
  XNOR2_X2 vscale_core_DW01_add_5_U337 ( .A(vscale_core_DW01_add_5n278), .B(vscale_core_DW01_add_5n40), .ZN(pipeline_md_N200) );
  NAND2_X2 vscale_core_DW01_add_5_U341 ( .A1(vscale_core_DW01_add_5n388), .A2(vscale_core_DW01_add_5n277), .ZN(vscale_core_DW01_add_5n40) );
  NAND2_X2 vscale_core_DW01_add_5_U344 ( .A1(pipeline_md_b[14]), .A2(pipeline_md_resp_result[14]), .ZN(vscale_core_DW01_add_5n277) );
  XOR2_X2 vscale_core_DW01_add_5_U345 ( .A(vscale_core_DW01_add_5n41), .B(vscale_core_DW01_add_5n285), .Z(pipeline_md_N199) );
  NAND2_X2 vscale_core_DW01_add_5_U351 ( .A1(vscale_core_DW01_add_5n389), .A2(vscale_core_DW01_add_5n284), .ZN(vscale_core_DW01_add_5n41) );
  NAND2_X2 vscale_core_DW01_add_5_U354 ( .A1(pipeline_md_b[13]), .A2(pipeline_md_resp_result[13]), .ZN(vscale_core_DW01_add_5n284) );
  XOR2_X2 vscale_core_DW01_add_5_U355 ( .A(vscale_core_DW01_add_5n42), .B(vscale_core_DW01_add_5n290), .Z(pipeline_md_N198) );
  NAND2_X2 vscale_core_DW01_add_5_U359 ( .A1(vscale_core_DW01_add_5n390), .A2(vscale_core_DW01_add_5n289), .ZN(vscale_core_DW01_add_5n42) );
  NAND2_X2 vscale_core_DW01_add_5_U362 ( .A1(pipeline_md_b[12]), .A2(pipeline_md_resp_result[12]), .ZN(vscale_core_DW01_add_5n289) );
  XOR2_X2 vscale_core_DW01_add_5_U363 ( .A(vscale_core_DW01_add_5n43), .B(vscale_core_DW01_add_5n298), .Z(pipeline_md_N197) );
  NAND2_X2 vscale_core_DW01_add_5_U366 ( .A1(vscale_core_DW01_add_5n306), .A2(vscale_core_DW01_add_5n294), .ZN(vscale_core_DW01_add_5n292) );
  NAND2_X2 vscale_core_DW01_add_5_U370 ( .A1(vscale_core_DW01_add_5n391), .A2(vscale_core_DW01_add_5n297), .ZN(vscale_core_DW01_add_5n43) );
  NAND2_X2 vscale_core_DW01_add_5_U373 ( .A1(pipeline_md_b[11]), .A2(pipeline_md_resp_result[11]), .ZN(vscale_core_DW01_add_5n297) );
  XNOR2_X2 vscale_core_DW01_add_5_U374 ( .A(vscale_core_DW01_add_5n303), .B(vscale_core_DW01_add_5n44), .ZN(pipeline_md_N196) );
  NAND2_X2 vscale_core_DW01_add_5_U378 ( .A1(vscale_core_DW01_add_5n392), .A2(vscale_core_DW01_add_5n302), .ZN(vscale_core_DW01_add_5n44) );
  NAND2_X2 vscale_core_DW01_add_5_U381 ( .A1(pipeline_md_b[10]), .A2(pipeline_md_resp_result[10]), .ZN(vscale_core_DW01_add_5n302) );
  XNOR2_X2 vscale_core_DW01_add_5_U382 ( .A(vscale_core_DW01_add_5n310), .B(vscale_core_DW01_add_5n45), .ZN(pipeline_md_N195) );
  NAND2_X2 vscale_core_DW01_add_5_U388 ( .A1(vscale_core_DW01_add_5n393), .A2(vscale_core_DW01_add_5n309), .ZN(vscale_core_DW01_add_5n45) );
  NAND2_X2 vscale_core_DW01_add_5_U391 ( .A1(pipeline_md_b[9]), .A2(pipeline_md_resp_result[9]), .ZN(vscale_core_DW01_add_5n309) );
  XOR2_X2 vscale_core_DW01_add_5_U392 ( .A(vscale_core_DW01_add_5n46), .B(vscale_core_DW01_add_5n313), .Z(pipeline_md_N194) );
  NAND2_X2 vscale_core_DW01_add_5_U394 ( .A1(vscale_core_DW01_add_5n394), .A2(vscale_core_DW01_add_5n312), .ZN(vscale_core_DW01_add_5n46) );
  NAND2_X2 vscale_core_DW01_add_5_U397 ( .A1(pipeline_md_b[8]), .A2(pipeline_md_resp_result[8]), .ZN(vscale_core_DW01_add_5n312) );
  XNOR2_X2 vscale_core_DW01_add_5_U398 ( .A(vscale_core_DW01_add_5n321), .B(vscale_core_DW01_add_5n47), .ZN(pipeline_md_N193) );
  NAND2_X2 vscale_core_DW01_add_5_U401 ( .A1(vscale_core_DW01_add_5n325), .A2(vscale_core_DW01_add_5n317), .ZN(vscale_core_DW01_add_5n315) );
  NAND2_X2 vscale_core_DW01_add_5_U405 ( .A1(vscale_core_DW01_add_5n395), .A2(vscale_core_DW01_add_5n320), .ZN(vscale_core_DW01_add_5n47) );
  NAND2_X2 vscale_core_DW01_add_5_U408 ( .A1(pipeline_md_b[7]), .A2(pipeline_md_resp_result[7]), .ZN(vscale_core_DW01_add_5n320) );
  XOR2_X2 vscale_core_DW01_add_5_U409 ( .A(vscale_core_DW01_add_5n48), .B(vscale_core_DW01_add_5n324), .Z(pipeline_md_N192) );
  NAND2_X2 vscale_core_DW01_add_5_U411 ( .A1(vscale_core_DW01_add_5n396), .A2(vscale_core_DW01_add_5n323), .ZN(vscale_core_DW01_add_5n48) );
  NAND2_X2 vscale_core_DW01_add_5_U414 ( .A1(pipeline_md_b[6]), .A2(pipeline_md_resp_result[6]), .ZN(vscale_core_DW01_add_5n323) );
  XOR2_X2 vscale_core_DW01_add_5_U415 ( .A(vscale_core_DW01_add_5n49), .B(vscale_core_DW01_add_5n329), .Z(pipeline_md_N191) );
  NAND2_X2 vscale_core_DW01_add_5_U419 ( .A1(vscale_core_DW01_add_5n397), .A2(vscale_core_DW01_add_5n328), .ZN(vscale_core_DW01_add_5n49) );
  NAND2_X2 vscale_core_DW01_add_5_U422 ( .A1(pipeline_md_b[5]), .A2(pipeline_md_resp_result[5]), .ZN(vscale_core_DW01_add_5n328) );
  XNOR2_X2 vscale_core_DW01_add_5_U423 ( .A(vscale_core_DW01_add_5n334), .B(vscale_core_DW01_add_5n50), .ZN(pipeline_md_N190) );
  NAND2_X2 vscale_core_DW01_add_5_U427 ( .A1(vscale_core_DW01_add_5n398), .A2(vscale_core_DW01_add_5n333), .ZN(vscale_core_DW01_add_5n50) );
  NAND2_X2 vscale_core_DW01_add_5_U430 ( .A1(pipeline_md_b[4]), .A2(pipeline_md_resp_result[4]), .ZN(vscale_core_DW01_add_5n333) );
  XNOR2_X2 vscale_core_DW01_add_5_U431 ( .A(vscale_core_DW01_add_5n340), .B(vscale_core_DW01_add_5n51), .ZN(pipeline_md_N189) );
  NAND2_X2 vscale_core_DW01_add_5_U436 ( .A1(vscale_core_DW01_add_5n399), .A2(vscale_core_DW01_add_5n339), .ZN(vscale_core_DW01_add_5n51) );
  NAND2_X2 vscale_core_DW01_add_5_U439 ( .A1(pipeline_md_b[3]), .A2(pipeline_md_resp_result[3]), .ZN(vscale_core_DW01_add_5n339) );
  XOR2_X2 vscale_core_DW01_add_5_U440 ( .A(vscale_core_DW01_add_5n52), .B(vscale_core_DW01_add_5n343), .Z(pipeline_md_N188) );
  NAND2_X2 vscale_core_DW01_add_5_U442 ( .A1(vscale_core_DW01_add_5n400), .A2(vscale_core_DW01_add_5n342), .ZN(vscale_core_DW01_add_5n52) );
  NAND2_X2 vscale_core_DW01_add_5_U445 ( .A1(pipeline_md_b[2]), .A2(pipeline_md_resp_result[2]), .ZN(vscale_core_DW01_add_5n342) );
  XOR2_X2 vscale_core_DW01_add_5_U446 ( .A(vscale_core_DW01_add_5n348), .B(vscale_core_DW01_add_5n53), .Z(pipeline_md_N187) );
  NAND2_X2 vscale_core_DW01_add_5_U449 ( .A1(vscale_core_DW01_add_5n401), .A2(vscale_core_DW01_add_5n346), .ZN(vscale_core_DW01_add_5n53) );
  NAND2_X2 vscale_core_DW01_add_5_U452 ( .A1(pipeline_md_b[1]), .A2(pipeline_md_resp_result[1]), .ZN(vscale_core_DW01_add_5n346) );
  NAND2_X2 vscale_core_DW01_add_5_U457 ( .A1(pipeline_md_b[0]), .A2(pipeline_md_resp_result[0]), .ZN(vscale_core_DW01_add_5n348) );
  AND2_X4 vscale_core_DW01_add_5_U461 ( .A1(vscale_core_DW01_add_5n607), .A2(vscale_core_DW01_add_5n348), .ZN(pipeline_md_N186) );
  NOR2_X2 vscale_core_DW01_add_5_U462 ( .A1(vscale_core_DW01_add_5n244), .A2(vscale_core_DW01_add_5n223), .ZN(vscale_core_DW01_add_5n221) );
  NOR2_X2 vscale_core_DW01_add_5_U463 ( .A1(vscale_core_DW01_add_5n154), .A2(vscale_core_DW01_add_5n129), .ZN(vscale_core_DW01_add_5n127) );
  AOI21_X2 vscale_core_DW01_add_5_U464 ( .B1(vscale_core_DW01_add_5n314), .B2(vscale_core_DW01_add_5n265), .A(vscale_core_DW01_add_5n266), .ZN(vscale_core_DW01_add_5n264) );
  NOR2_X2 vscale_core_DW01_add_5_U465 ( .A1(vscale_core_DW01_add_5n292), .A2(vscale_core_DW01_add_5n267), .ZN(vscale_core_DW01_add_5n265) );
  OAI21_X2 vscale_core_DW01_add_5_U466 ( .B1(vscale_core_DW01_add_5n293), .B2(vscale_core_DW01_add_5n267), .A(vscale_core_DW01_add_5n268), .ZN(vscale_core_DW01_add_5n266) );
  OAI21_X2 vscale_core_DW01_add_5_U467 ( .B1(vscale_core_DW01_add_5n264), .B2(vscale_core_DW01_add_5n177), .A(vscale_core_DW01_add_5n178), .ZN(vscale_core_DW01_add_5n176) );
  AOI21_X2 vscale_core_DW01_add_5_U468 ( .B1(vscale_core_DW01_add_5n222), .B2(vscale_core_DW01_add_5n179), .A(vscale_core_DW01_add_5n180), .ZN(vscale_core_DW01_add_5n178) );
  NOR2_X2 vscale_core_DW01_add_5_U469 ( .A1(vscale_core_DW01_add_5n202), .A2(vscale_core_DW01_add_5n181), .ZN(vscale_core_DW01_add_5n179) );
  AOI21_X2 vscale_core_DW01_add_5_U470 ( .B1(vscale_core_DW01_add_5n219), .B2(vscale_core_DW01_add_5n212), .A(vscale_core_DW01_add_5n213), .ZN(vscale_core_DW01_add_5n211) );
  AOI21_X2 vscale_core_DW01_add_5_U471 ( .B1(vscale_core_DW01_add_5n240), .B2(vscale_core_DW01_add_5n233), .A(vscale_core_DW01_add_5n234), .ZN(vscale_core_DW01_add_5n232) );
  AOI21_X2 vscale_core_DW01_add_5_U472 ( .B1(vscale_core_DW01_add_5n263), .B2(vscale_core_DW01_add_5n254), .A(vscale_core_DW01_add_5n255), .ZN(vscale_core_DW01_add_5n253) );
  AOI21_X2 vscale_core_DW01_add_5_U473 ( .B1(vscale_core_DW01_add_5n198), .B2(vscale_core_DW01_add_5n191), .A(vscale_core_DW01_add_5n192), .ZN(vscale_core_DW01_add_5n190) );
  AOI21_X2 vscale_core_DW01_add_5_U474 ( .B1(vscale_core_DW01_add_5n263), .B2(vscale_core_DW01_add_5n242), .A(vscale_core_DW01_add_5n243), .ZN(vscale_core_DW01_add_5n241) );
  AOI21_X2 vscale_core_DW01_add_5_U475 ( .B1(vscale_core_DW01_add_5n219), .B2(vscale_core_DW01_add_5n200), .A(vscale_core_DW01_add_5n201), .ZN(vscale_core_DW01_add_5n199) );
  AOI21_X2 vscale_core_DW01_add_5_U476 ( .B1(vscale_core_DW01_add_5n263), .B2(vscale_core_DW01_add_5n221), .A(vscale_core_DW01_add_5n222), .ZN(vscale_core_DW01_add_5n220) );
  OAI21_X2 vscale_core_DW01_add_5_U477 ( .B1(vscale_core_DW01_add_5n313), .B2(vscale_core_DW01_add_5n292), .A(vscale_core_DW01_add_5n293), .ZN(vscale_core_DW01_add_5n291) );
  OAI21_X2 vscale_core_DW01_add_5_U478 ( .B1(vscale_core_DW01_add_5n175), .B2(vscale_core_DW01_add_5n154), .A(vscale_core_DW01_add_5n155), .ZN(vscale_core_DW01_add_5n153) );
  OAI21_X2 vscale_core_DW01_add_5_U479 ( .B1(vscale_core_DW01_add_5n290), .B2(vscale_core_DW01_add_5n279), .A(vscale_core_DW01_add_5n280), .ZN(vscale_core_DW01_add_5n278) );
  OAI21_X2 vscale_core_DW01_add_5_U480 ( .B1(vscale_core_DW01_add_5n313), .B2(vscale_core_DW01_add_5n304), .A(vscale_core_DW01_add_5n305), .ZN(vscale_core_DW01_add_5n303) );
  OAI21_X2 vscale_core_DW01_add_5_U481 ( .B1(vscale_core_DW01_add_5n175), .B2(vscale_core_DW01_add_5n125), .A(vscale_core_DW01_add_5n126), .ZN(vscale_core_DW01_add_5n124) );
  OAI21_X2 vscale_core_DW01_add_5_U482 ( .B1(vscale_core_DW01_add_5n152), .B2(vscale_core_DW01_add_5n141), .A(vscale_core_DW01_add_5n142), .ZN(vscale_core_DW01_add_5n140) );
  OAI21_X2 vscale_core_DW01_add_5_U483 ( .B1(vscale_core_DW01_add_5n175), .B2(vscale_core_DW01_add_5n166), .A(vscale_core_DW01_add_5n167), .ZN(vscale_core_DW01_add_5n165) );
  OAI21_X2 vscale_core_DW01_add_5_U484 ( .B1(vscale_core_DW01_add_5n175), .B2(vscale_core_DW01_add_5n113), .A(vscale_core_DW01_add_5n114), .ZN(vscale_core_DW01_add_5n112) );
  AOI21_X2 vscale_core_DW01_add_5_U485 ( .B1(vscale_core_DW01_add_5n334), .B2(vscale_core_DW01_add_5n325), .A(vscale_core_DW01_add_5n326), .ZN(vscale_core_DW01_add_5n324) );
  AOI21_X2 vscale_core_DW01_add_5_U486 ( .B1(vscale_core_DW01_add_5n72), .B2(vscale_core_DW01_add_5n606), .A(vscale_core_DW01_add_5n69), .ZN(vscale_core_DW01_add_5n67) );
  AOI21_X2 vscale_core_DW01_add_5_U487 ( .B1(vscale_core_DW01_add_5n80), .B2(vscale_core_DW01_add_5n603), .A(vscale_core_DW01_add_5n77), .ZN(vscale_core_DW01_add_5n75) );
  AOI21_X2 vscale_core_DW01_add_5_U488 ( .B1(vscale_core_DW01_add_5n88), .B2(vscale_core_DW01_add_5n605), .A(vscale_core_DW01_add_5n85), .ZN(vscale_core_DW01_add_5n83) );
  AOI21_X2 vscale_core_DW01_add_5_U489 ( .B1(vscale_core_DW01_add_5n96), .B2(vscale_core_DW01_add_5n604), .A(vscale_core_DW01_add_5n93), .ZN(vscale_core_DW01_add_5n91) );
  AOI21_X2 vscale_core_DW01_add_5_U490 ( .B1(vscale_core_DW01_add_5n104), .B2(vscale_core_DW01_add_5n602), .A(vscale_core_DW01_add_5n101), .ZN(vscale_core_DW01_add_5n99) );
  AOI21_X2 vscale_core_DW01_add_5_U491 ( .B1(vscale_core_DW01_add_5n176), .B2(vscale_core_DW01_add_5n108), .A(vscale_core_DW01_add_5n109), .ZN(vscale_core_DW01_add_5n107) );
  NOR2_X2 vscale_core_DW01_add_5_U492 ( .A1(vscale_core_DW01_add_5n113), .A2(vscale_core_DW01_add_5n110), .ZN(vscale_core_DW01_add_5n108) );
  OAI21_X2 vscale_core_DW01_add_5_U493 ( .B1(vscale_core_DW01_add_5n114), .B2(vscale_core_DW01_add_5n110), .A(vscale_core_DW01_add_5n111), .ZN(vscale_core_DW01_add_5n109) );
  AOI21_X2 vscale_core_DW01_add_5_U494 ( .B1(vscale_core_DW01_add_5n156), .B2(vscale_core_DW01_add_5n169), .A(vscale_core_DW01_add_5n157), .ZN(vscale_core_DW01_add_5n155) );
  OAI21_X2 vscale_core_DW01_add_5_U495 ( .B1(vscale_core_DW01_add_5n158), .B2(vscale_core_DW01_add_5n164), .A(vscale_core_DW01_add_5n159), .ZN(vscale_core_DW01_add_5n157) );
  AOI21_X2 vscale_core_DW01_add_5_U496 ( .B1(vscale_core_DW01_add_5n294), .B2(vscale_core_DW01_add_5n307), .A(vscale_core_DW01_add_5n295), .ZN(vscale_core_DW01_add_5n293) );
  OAI21_X2 vscale_core_DW01_add_5_U497 ( .B1(vscale_core_DW01_add_5n296), .B2(vscale_core_DW01_add_5n302), .A(vscale_core_DW01_add_5n297), .ZN(vscale_core_DW01_add_5n295) );
  AOI21_X2 vscale_core_DW01_add_5_U498 ( .B1(vscale_core_DW01_add_5n128), .B2(vscale_core_DW01_add_5n115), .A(vscale_core_DW01_add_5n116), .ZN(vscale_core_DW01_add_5n114) );
  OAI21_X2 vscale_core_DW01_add_5_U499 ( .B1(vscale_core_DW01_add_5n117), .B2(vscale_core_DW01_add_5n123), .A(vscale_core_DW01_add_5n118), .ZN(vscale_core_DW01_add_5n116) );
  AOI21_X2 vscale_core_DW01_add_5_U500 ( .B1(vscale_core_DW01_add_5n336), .B2(vscale_core_DW01_add_5n344), .A(vscale_core_DW01_add_5n337), .ZN(vscale_core_DW01_add_5n335) );
  NOR2_X2 vscale_core_DW01_add_5_U501 ( .A1(vscale_core_DW01_add_5n341), .A2(vscale_core_DW01_add_5n338), .ZN(vscale_core_DW01_add_5n336) );
  OAI21_X2 vscale_core_DW01_add_5_U502 ( .B1(vscale_core_DW01_add_5n338), .B2(vscale_core_DW01_add_5n342), .A(vscale_core_DW01_add_5n339), .ZN(vscale_core_DW01_add_5n337) );
  AOI21_X2 vscale_core_DW01_add_5_U503 ( .B1(vscale_core_DW01_add_5n204), .B2(vscale_core_DW01_add_5n213), .A(vscale_core_DW01_add_5n205), .ZN(vscale_core_DW01_add_5n203) );
  OAI21_X2 vscale_core_DW01_add_5_U504 ( .B1(vscale_core_DW01_add_5n206), .B2(vscale_core_DW01_add_5n210), .A(vscale_core_DW01_add_5n207), .ZN(vscale_core_DW01_add_5n205) );
  AOI21_X2 vscale_core_DW01_add_5_U505 ( .B1(vscale_core_DW01_add_5n246), .B2(vscale_core_DW01_add_5n255), .A(vscale_core_DW01_add_5n247), .ZN(vscale_core_DW01_add_5n245) );
  OAI21_X2 vscale_core_DW01_add_5_U506 ( .B1(vscale_core_DW01_add_5n248), .B2(vscale_core_DW01_add_5n252), .A(vscale_core_DW01_add_5n249), .ZN(vscale_core_DW01_add_5n247) );
  OAI21_X2 vscale_core_DW01_add_5_U507 ( .B1(vscale_core_DW01_add_5n245), .B2(vscale_core_DW01_add_5n223), .A(vscale_core_DW01_add_5n224), .ZN(vscale_core_DW01_add_5n222) );
  AOI21_X2 vscale_core_DW01_add_5_U508 ( .B1(vscale_core_DW01_add_5n225), .B2(vscale_core_DW01_add_5n234), .A(vscale_core_DW01_add_5n226), .ZN(vscale_core_DW01_add_5n224) );
  OAI21_X2 vscale_core_DW01_add_5_U509 ( .B1(vscale_core_DW01_add_5n227), .B2(vscale_core_DW01_add_5n231), .A(vscale_core_DW01_add_5n228), .ZN(vscale_core_DW01_add_5n226) );
  OAI21_X2 vscale_core_DW01_add_5_U510 ( .B1(vscale_core_DW01_add_5n155), .B2(vscale_core_DW01_add_5n129), .A(vscale_core_DW01_add_5n130), .ZN(vscale_core_DW01_add_5n128) );
  AOI21_X2 vscale_core_DW01_add_5_U511 ( .B1(vscale_core_DW01_add_5n131), .B2(vscale_core_DW01_add_5n144), .A(vscale_core_DW01_add_5n132), .ZN(vscale_core_DW01_add_5n130) );
  OAI21_X2 vscale_core_DW01_add_5_U512 ( .B1(vscale_core_DW01_add_5n133), .B2(vscale_core_DW01_add_5n139), .A(vscale_core_DW01_add_5n134), .ZN(vscale_core_DW01_add_5n132) );
  OAI21_X2 vscale_core_DW01_add_5_U513 ( .B1(vscale_core_DW01_add_5n335), .B2(vscale_core_DW01_add_5n315), .A(vscale_core_DW01_add_5n316), .ZN(vscale_core_DW01_add_5n314) );
  AOI21_X2 vscale_core_DW01_add_5_U514 ( .B1(vscale_core_DW01_add_5n317), .B2(vscale_core_DW01_add_5n326), .A(vscale_core_DW01_add_5n318), .ZN(vscale_core_DW01_add_5n316) );
  NOR2_X2 vscale_core_DW01_add_5_U515 ( .A1(vscale_core_DW01_add_5n322), .A2(vscale_core_DW01_add_5n319), .ZN(vscale_core_DW01_add_5n317) );
  OAI21_X2 vscale_core_DW01_add_5_U516 ( .B1(vscale_core_DW01_add_5n75), .B2(vscale_core_DW01_add_5n73), .A(vscale_core_DW01_add_5n74), .ZN(vscale_core_DW01_add_5n72) );
  OAI21_X2 vscale_core_DW01_add_5_U517 ( .B1(vscale_core_DW01_add_5n83), .B2(vscale_core_DW01_add_5n81), .A(vscale_core_DW01_add_5n82), .ZN(vscale_core_DW01_add_5n80) );
  OAI21_X2 vscale_core_DW01_add_5_U518 ( .B1(vscale_core_DW01_add_5n91), .B2(vscale_core_DW01_add_5n89), .A(vscale_core_DW01_add_5n90), .ZN(vscale_core_DW01_add_5n88) );
  OAI21_X2 vscale_core_DW01_add_5_U519 ( .B1(vscale_core_DW01_add_5n99), .B2(vscale_core_DW01_add_5n97), .A(vscale_core_DW01_add_5n98), .ZN(vscale_core_DW01_add_5n96) );
  OAI21_X2 vscale_core_DW01_add_5_U520 ( .B1(vscale_core_DW01_add_5n107), .B2(vscale_core_DW01_add_5n105), .A(vscale_core_DW01_add_5n106), .ZN(vscale_core_DW01_add_5n104) );
  OAI21_X2 vscale_core_DW01_add_5_U521 ( .B1(vscale_core_DW01_add_5n327), .B2(vscale_core_DW01_add_5n333), .A(vscale_core_DW01_add_5n328), .ZN(vscale_core_DW01_add_5n326) );
  OAI21_X2 vscale_core_DW01_add_5_U522 ( .B1(vscale_core_DW01_add_5n214), .B2(vscale_core_DW01_add_5n218), .A(vscale_core_DW01_add_5n215), .ZN(vscale_core_DW01_add_5n213) );
  OAI21_X2 vscale_core_DW01_add_5_U523 ( .B1(vscale_core_DW01_add_5n193), .B2(vscale_core_DW01_add_5n197), .A(vscale_core_DW01_add_5n194), .ZN(vscale_core_DW01_add_5n192) );
  OAI21_X2 vscale_core_DW01_add_5_U524 ( .B1(vscale_core_DW01_add_5n235), .B2(vscale_core_DW01_add_5n239), .A(vscale_core_DW01_add_5n236), .ZN(vscale_core_DW01_add_5n234) );
  OAI21_X2 vscale_core_DW01_add_5_U525 ( .B1(vscale_core_DW01_add_5n256), .B2(vscale_core_DW01_add_5n262), .A(vscale_core_DW01_add_5n257), .ZN(vscale_core_DW01_add_5n255) );
  OAI21_X2 vscale_core_DW01_add_5_U526 ( .B1(vscale_core_DW01_add_5n170), .B2(vscale_core_DW01_add_5n174), .A(vscale_core_DW01_add_5n171), .ZN(vscale_core_DW01_add_5n169) );
  OAI21_X2 vscale_core_DW01_add_5_U527 ( .B1(vscale_core_DW01_add_5n145), .B2(vscale_core_DW01_add_5n151), .A(vscale_core_DW01_add_5n146), .ZN(vscale_core_DW01_add_5n144) );
  OAI21_X2 vscale_core_DW01_add_5_U528 ( .B1(vscale_core_DW01_add_5n308), .B2(vscale_core_DW01_add_5n312), .A(vscale_core_DW01_add_5n309), .ZN(vscale_core_DW01_add_5n307) );
  OAI21_X2 vscale_core_DW01_add_5_U529 ( .B1(vscale_core_DW01_add_5n283), .B2(vscale_core_DW01_add_5n289), .A(vscale_core_DW01_add_5n284), .ZN(vscale_core_DW01_add_5n282) );
  OAI21_X2 vscale_core_DW01_add_5_U530 ( .B1(vscale_core_DW01_add_5n345), .B2(vscale_core_DW01_add_5n348), .A(vscale_core_DW01_add_5n346), .ZN(vscale_core_DW01_add_5n344) );
  AOI21_X2 vscale_core_DW01_add_5_U531 ( .B1(vscale_core_DW01_add_5n269), .B2(vscale_core_DW01_add_5n282), .A(vscale_core_DW01_add_5n270), .ZN(vscale_core_DW01_add_5n268) );
  OAI21_X2 vscale_core_DW01_add_5_U532 ( .B1(vscale_core_DW01_add_5n271), .B2(vscale_core_DW01_add_5n277), .A(vscale_core_DW01_add_5n272), .ZN(vscale_core_DW01_add_5n270) );
  OAI21_X2 vscale_core_DW01_add_5_U533 ( .B1(vscale_core_DW01_add_5n319), .B2(vscale_core_DW01_add_5n323), .A(vscale_core_DW01_add_5n320), .ZN(vscale_core_DW01_add_5n318) );
  OAI21_X2 vscale_core_DW01_add_5_U534 ( .B1(vscale_core_DW01_add_5n203), .B2(vscale_core_DW01_add_5n181), .A(vscale_core_DW01_add_5n182), .ZN(vscale_core_DW01_add_5n180) );
  AOI21_X2 vscale_core_DW01_add_5_U535 ( .B1(vscale_core_DW01_add_5n183), .B2(vscale_core_DW01_add_5n192), .A(vscale_core_DW01_add_5n184), .ZN(vscale_core_DW01_add_5n182) );
  OAI21_X2 vscale_core_DW01_add_5_U536 ( .B1(vscale_core_DW01_add_5n185), .B2(vscale_core_DW01_add_5n189), .A(vscale_core_DW01_add_5n186), .ZN(vscale_core_DW01_add_5n184) );
  NOR2_X2 vscale_core_DW01_add_5_U537 ( .A1(vscale_core_DW01_add_5n276), .A2(vscale_core_DW01_add_5n271), .ZN(vscale_core_DW01_add_5n269) );
  NOR2_X2 vscale_core_DW01_add_5_U538 ( .A1(vscale_core_DW01_add_5n301), .A2(vscale_core_DW01_add_5n296), .ZN(vscale_core_DW01_add_5n294) );
  NOR2_X2 vscale_core_DW01_add_5_U539 ( .A1(vscale_core_DW01_add_5n188), .A2(vscale_core_DW01_add_5n185), .ZN(vscale_core_DW01_add_5n183) );
  NOR2_X2 vscale_core_DW01_add_5_U540 ( .A1(vscale_core_DW01_add_5n209), .A2(vscale_core_DW01_add_5n206), .ZN(vscale_core_DW01_add_5n204) );
  NOR2_X2 vscale_core_DW01_add_5_U541 ( .A1(vscale_core_DW01_add_5n230), .A2(vscale_core_DW01_add_5n227), .ZN(vscale_core_DW01_add_5n225) );
  NOR2_X2 vscale_core_DW01_add_5_U542 ( .A1(vscale_core_DW01_add_5n251), .A2(vscale_core_DW01_add_5n248), .ZN(vscale_core_DW01_add_5n246) );
  NOR2_X2 vscale_core_DW01_add_5_U543 ( .A1(vscale_core_DW01_add_5n138), .A2(vscale_core_DW01_add_5n133), .ZN(vscale_core_DW01_add_5n131) );
  NOR2_X2 vscale_core_DW01_add_5_U544 ( .A1(vscale_core_DW01_add_5n163), .A2(vscale_core_DW01_add_5n158), .ZN(vscale_core_DW01_add_5n156) );
  NOR2_X2 vscale_core_DW01_add_5_U545 ( .A1(vscale_core_DW01_add_5n196), .A2(vscale_core_DW01_add_5n193), .ZN(vscale_core_DW01_add_5n191) );
  NOR2_X2 vscale_core_DW01_add_5_U546 ( .A1(vscale_core_DW01_add_5n217), .A2(vscale_core_DW01_add_5n214), .ZN(vscale_core_DW01_add_5n212) );
  NOR2_X2 vscale_core_DW01_add_5_U547 ( .A1(vscale_core_DW01_add_5n238), .A2(vscale_core_DW01_add_5n235), .ZN(vscale_core_DW01_add_5n233) );
  NOR2_X2 vscale_core_DW01_add_5_U548 ( .A1(vscale_core_DW01_add_5n288), .A2(vscale_core_DW01_add_5n283), .ZN(vscale_core_DW01_add_5n281) );
  NOR2_X2 vscale_core_DW01_add_5_U549 ( .A1(vscale_core_DW01_add_5n311), .A2(vscale_core_DW01_add_5n308), .ZN(vscale_core_DW01_add_5n306) );
  NOR2_X2 vscale_core_DW01_add_5_U550 ( .A1(vscale_core_DW01_add_5n150), .A2(vscale_core_DW01_add_5n145), .ZN(vscale_core_DW01_add_5n143) );
  NOR2_X2 vscale_core_DW01_add_5_U551 ( .A1(vscale_core_DW01_add_5n332), .A2(vscale_core_DW01_add_5n327), .ZN(vscale_core_DW01_add_5n325) );
  NOR2_X2 vscale_core_DW01_add_5_U552 ( .A1(vscale_core_DW01_add_5n261), .A2(vscale_core_DW01_add_5n256), .ZN(vscale_core_DW01_add_5n254) );
  NOR2_X2 vscale_core_DW01_add_5_U553 ( .A1(vscale_core_DW01_add_5n122), .A2(vscale_core_DW01_add_5n117), .ZN(vscale_core_DW01_add_5n115) );
  NOR2_X2 vscale_core_DW01_add_5_U554 ( .A1(vscale_core_DW01_add_5n173), .A2(vscale_core_DW01_add_5n170), .ZN(vscale_core_DW01_add_5n168) );
  AOI21_X2 vscale_core_DW01_add_5_U555 ( .B1(vscale_core_DW01_add_5n124), .B2(vscale_core_DW01_add_5n362), .A(vscale_core_DW01_add_5n121), .ZN(vscale_core_DW01_add_5n119) );
  AOI21_X2 vscale_core_DW01_add_5_U556 ( .B1(vscale_core_DW01_add_5n140), .B2(vscale_core_DW01_add_5n364), .A(vscale_core_DW01_add_5n137), .ZN(vscale_core_DW01_add_5n135) );
  AOI21_X2 vscale_core_DW01_add_5_U557 ( .B1(vscale_core_DW01_add_5n153), .B2(vscale_core_DW01_add_5n366), .A(vscale_core_DW01_add_5n149), .ZN(vscale_core_DW01_add_5n147) );
  AOI21_X2 vscale_core_DW01_add_5_U558 ( .B1(vscale_core_DW01_add_5n165), .B2(vscale_core_DW01_add_5n368), .A(vscale_core_DW01_add_5n162), .ZN(vscale_core_DW01_add_5n160) );
  AOI21_X2 vscale_core_DW01_add_5_U559 ( .B1(vscale_core_DW01_add_5n263), .B2(vscale_core_DW01_add_5n386), .A(vscale_core_DW01_add_5n260), .ZN(vscale_core_DW01_add_5n258) );
  AOI21_X2 vscale_core_DW01_add_5_U560 ( .B1(vscale_core_DW01_add_5n278), .B2(vscale_core_DW01_add_5n388), .A(vscale_core_DW01_add_5n275), .ZN(vscale_core_DW01_add_5n273) );
  AOI21_X2 vscale_core_DW01_add_5_U561 ( .B1(vscale_core_DW01_add_5n291), .B2(vscale_core_DW01_add_5n390), .A(vscale_core_DW01_add_5n287), .ZN(vscale_core_DW01_add_5n285) );
  AOI21_X2 vscale_core_DW01_add_5_U562 ( .B1(vscale_core_DW01_add_5n303), .B2(vscale_core_DW01_add_5n392), .A(vscale_core_DW01_add_5n300), .ZN(vscale_core_DW01_add_5n298) );
  OAI21_X2 vscale_core_DW01_add_5_U563 ( .B1(vscale_core_DW01_add_5n211), .B2(vscale_core_DW01_add_5n209), .A(vscale_core_DW01_add_5n210), .ZN(vscale_core_DW01_add_5n208) );
  OAI21_X2 vscale_core_DW01_add_5_U564 ( .B1(vscale_core_DW01_add_5n220), .B2(vscale_core_DW01_add_5n217), .A(vscale_core_DW01_add_5n218), .ZN(vscale_core_DW01_add_5n216) );
  OAI21_X2 vscale_core_DW01_add_5_U565 ( .B1(vscale_core_DW01_add_5n232), .B2(vscale_core_DW01_add_5n230), .A(vscale_core_DW01_add_5n231), .ZN(vscale_core_DW01_add_5n229) );
  OAI21_X2 vscale_core_DW01_add_5_U566 ( .B1(vscale_core_DW01_add_5n241), .B2(vscale_core_DW01_add_5n238), .A(vscale_core_DW01_add_5n239), .ZN(vscale_core_DW01_add_5n237) );
  OAI21_X2 vscale_core_DW01_add_5_U567 ( .B1(vscale_core_DW01_add_5n253), .B2(vscale_core_DW01_add_5n251), .A(vscale_core_DW01_add_5n252), .ZN(vscale_core_DW01_add_5n250) );
  OAI21_X2 vscale_core_DW01_add_5_U568 ( .B1(vscale_core_DW01_add_5n199), .B2(vscale_core_DW01_add_5n196), .A(vscale_core_DW01_add_5n197), .ZN(vscale_core_DW01_add_5n195) );
  OAI21_X2 vscale_core_DW01_add_5_U569 ( .B1(vscale_core_DW01_add_5n190), .B2(vscale_core_DW01_add_5n188), .A(vscale_core_DW01_add_5n189), .ZN(vscale_core_DW01_add_5n187) );
  OAI21_X2 vscale_core_DW01_add_5_U570 ( .B1(vscale_core_DW01_add_5n175), .B2(vscale_core_DW01_add_5n173), .A(vscale_core_DW01_add_5n174), .ZN(vscale_core_DW01_add_5n172) );
  AOI21_X2 vscale_core_DW01_add_5_U571 ( .B1(vscale_core_DW01_add_5n334), .B2(vscale_core_DW01_add_5n398), .A(vscale_core_DW01_add_5n331), .ZN(vscale_core_DW01_add_5n329) );
  OAI21_X2 vscale_core_DW01_add_5_U572 ( .B1(vscale_core_DW01_add_5n324), .B2(vscale_core_DW01_add_5n322), .A(vscale_core_DW01_add_5n323), .ZN(vscale_core_DW01_add_5n321) );
  OAI21_X2 vscale_core_DW01_add_5_U573 ( .B1(vscale_core_DW01_add_5n343), .B2(vscale_core_DW01_add_5n341), .A(vscale_core_DW01_add_5n342), .ZN(vscale_core_DW01_add_5n340) );
  OAI21_X2 vscale_core_DW01_add_5_U574 ( .B1(vscale_core_DW01_add_5n313), .B2(vscale_core_DW01_add_5n311), .A(vscale_core_DW01_add_5n312), .ZN(vscale_core_DW01_add_5n310) );
  NOR2_X2 vscale_core_DW01_add_5_U575 ( .A1(pipeline_md_b[39]), .A2(pipeline_md_result[39]), .ZN(vscale_core_DW01_add_5n133) );
  NOR2_X2 vscale_core_DW01_add_5_U576 ( .A1(pipeline_md_b[37]), .A2(pipeline_md_result[37]), .ZN(vscale_core_DW01_add_5n145) );
  NOR2_X2 vscale_core_DW01_add_5_U577 ( .A1(pipeline_md_b[35]), .A2(pipeline_md_result[35]), .ZN(vscale_core_DW01_add_5n158) );
  NOR2_X2 vscale_core_DW01_add_5_U578 ( .A1(pipeline_md_b[33]), .A2(pipeline_md_result[33]), .ZN(vscale_core_DW01_add_5n170) );
  NOR2_X2 vscale_core_DW01_add_5_U579 ( .A1(pipeline_md_b[27]), .A2(pipeline_md_resp_result[27]), .ZN(vscale_core_DW01_add_5n206) );
  NOR2_X2 vscale_core_DW01_add_5_U580 ( .A1(pipeline_md_b[25]), .A2(pipeline_md_resp_result[25]), .ZN(vscale_core_DW01_add_5n214) );
  NOR2_X2 vscale_core_DW01_add_5_U581 ( .A1(pipeline_md_b[23]), .A2(pipeline_md_resp_result[23]), .ZN(vscale_core_DW01_add_5n227) );
  NOR2_X2 vscale_core_DW01_add_5_U582 ( .A1(pipeline_md_b[21]), .A2(pipeline_md_resp_result[21]), .ZN(vscale_core_DW01_add_5n235) );
  NOR2_X2 vscale_core_DW01_add_5_U583 ( .A1(pipeline_md_b[19]), .A2(pipeline_md_resp_result[19]), .ZN(vscale_core_DW01_add_5n248) );
  NOR2_X2 vscale_core_DW01_add_5_U584 ( .A1(pipeline_md_b[17]), .A2(pipeline_md_resp_result[17]), .ZN(vscale_core_DW01_add_5n256) );
  NOR2_X2 vscale_core_DW01_add_5_U585 ( .A1(pipeline_md_b[15]), .A2(pipeline_md_resp_result[15]), .ZN(vscale_core_DW01_add_5n271) );
  NOR2_X2 vscale_core_DW01_add_5_U586 ( .A1(pipeline_md_b[13]), .A2(pipeline_md_resp_result[13]), .ZN(vscale_core_DW01_add_5n283) );
  NOR2_X2 vscale_core_DW01_add_5_U587 ( .A1(pipeline_md_b[11]), .A2(pipeline_md_resp_result[11]), .ZN(vscale_core_DW01_add_5n296) );
  NOR2_X2 vscale_core_DW01_add_5_U588 ( .A1(pipeline_md_b[9]), .A2(pipeline_md_resp_result[9]), .ZN(vscale_core_DW01_add_5n308) );
  NOR2_X2 vscale_core_DW01_add_5_U589 ( .A1(pipeline_md_b[7]), .A2(pipeline_md_resp_result[7]), .ZN(vscale_core_DW01_add_5n319) );
  NOR2_X2 vscale_core_DW01_add_5_U590 ( .A1(pipeline_md_b[5]), .A2(pipeline_md_resp_result[5]), .ZN(vscale_core_DW01_add_5n327) );
  NOR2_X2 vscale_core_DW01_add_5_U591 ( .A1(pipeline_md_b[3]), .A2(pipeline_md_resp_result[3]), .ZN(vscale_core_DW01_add_5n338) );
  NOR2_X2 vscale_core_DW01_add_5_U592 ( .A1(pipeline_md_b[29]), .A2(pipeline_md_resp_result[29]), .ZN(vscale_core_DW01_add_5n193) );
  NOR2_X2 vscale_core_DW01_add_5_U593 ( .A1(pipeline_md_b[31]), .A2(pipeline_md_resp_result[31]), .ZN(vscale_core_DW01_add_5n185) );
  OAI21_X2 vscale_core_DW01_add_5_U594 ( .B1(vscale_core_DW01_add_5n67), .B2(vscale_core_DW01_add_5n65), .A(vscale_core_DW01_add_5n66), .ZN(vscale_core_DW01_add_5n64) );
  NOR2_X2 vscale_core_DW01_add_5_U595 ( .A1(pipeline_md_b[26]), .A2(pipeline_md_resp_result[26]), .ZN(vscale_core_DW01_add_5n209) );
  NOR2_X2 vscale_core_DW01_add_5_U596 ( .A1(pipeline_md_b[22]), .A2(pipeline_md_resp_result[22]), .ZN(vscale_core_DW01_add_5n230) );
  NOR2_X2 vscale_core_DW01_add_5_U597 ( .A1(pipeline_md_b[20]), .A2(pipeline_md_resp_result[20]), .ZN(vscale_core_DW01_add_5n238) );
  NOR2_X2 vscale_core_DW01_add_5_U598 ( .A1(pipeline_md_b[18]), .A2(pipeline_md_resp_result[18]), .ZN(vscale_core_DW01_add_5n251) );
  NOR2_X2 vscale_core_DW01_add_5_U599 ( .A1(pipeline_md_b[8]), .A2(pipeline_md_resp_result[8]), .ZN(vscale_core_DW01_add_5n311) );
  NOR2_X2 vscale_core_DW01_add_5_U600 ( .A1(pipeline_md_b[6]), .A2(pipeline_md_resp_result[6]), .ZN(vscale_core_DW01_add_5n322) );
  NOR2_X2 vscale_core_DW01_add_5_U601 ( .A1(pipeline_md_b[2]), .A2(pipeline_md_resp_result[2]), .ZN(vscale_core_DW01_add_5n341) );
  NOR2_X2 vscale_core_DW01_add_5_U602 ( .A1(pipeline_md_b[28]), .A2(pipeline_md_resp_result[28]), .ZN(vscale_core_DW01_add_5n196) );
  NOR2_X2 vscale_core_DW01_add_5_U603 ( .A1(pipeline_md_b[30]), .A2(pipeline_md_resp_result[30]), .ZN(vscale_core_DW01_add_5n188) );
  NOR2_X2 vscale_core_DW01_add_5_U604 ( .A1(pipeline_md_b[1]), .A2(pipeline_md_resp_result[1]), .ZN(vscale_core_DW01_add_5n345) );
  NOR2_X2 vscale_core_DW01_add_5_U605 ( .A1(pipeline_md_b[14]), .A2(pipeline_md_resp_result[14]), .ZN(vscale_core_DW01_add_5n276) );
  NOR2_X2 vscale_core_DW01_add_5_U606 ( .A1(pipeline_md_b[12]), .A2(pipeline_md_resp_result[12]), .ZN(vscale_core_DW01_add_5n288) );
  NOR2_X2 vscale_core_DW01_add_5_U607 ( .A1(pipeline_md_b[10]), .A2(pipeline_md_resp_result[10]), .ZN(vscale_core_DW01_add_5n301) );
  NOR2_X2 vscale_core_DW01_add_5_U608 ( .A1(pipeline_md_b[38]), .A2(pipeline_md_result[38]), .ZN(vscale_core_DW01_add_5n138) );
  NOR2_X2 vscale_core_DW01_add_5_U609 ( .A1(pipeline_md_b[36]), .A2(pipeline_md_result[36]), .ZN(vscale_core_DW01_add_5n150) );
  NOR2_X2 vscale_core_DW01_add_5_U610 ( .A1(pipeline_md_b[34]), .A2(pipeline_md_result[34]), .ZN(vscale_core_DW01_add_5n163) );
  NOR2_X2 vscale_core_DW01_add_5_U611 ( .A1(pipeline_md_b[41]), .A2(pipeline_md_result[41]), .ZN(vscale_core_DW01_add_5n117) );
  NOR2_X2 vscale_core_DW01_add_5_U612 ( .A1(pipeline_md_b[32]), .A2(pipeline_md_result[32]), .ZN(vscale_core_DW01_add_5n173) );
  NOR2_X2 vscale_core_DW01_add_5_U613 ( .A1(pipeline_md_b[24]), .A2(pipeline_md_resp_result[24]), .ZN(vscale_core_DW01_add_5n217) );
  NOR2_X2 vscale_core_DW01_add_5_U614 ( .A1(pipeline_md_b[42]), .A2(pipeline_md_result[42]), .ZN(vscale_core_DW01_add_5n110) );
  NOR2_X2 vscale_core_DW01_add_5_U615 ( .A1(pipeline_md_b[4]), .A2(pipeline_md_resp_result[4]), .ZN(vscale_core_DW01_add_5n332) );
  NOR2_X2 vscale_core_DW01_add_5_U616 ( .A1(pipeline_md_b[16]), .A2(pipeline_md_resp_result[16]), .ZN(vscale_core_DW01_add_5n261) );
  NOR2_X2 vscale_core_DW01_add_5_U617 ( .A1(pipeline_md_b[40]), .A2(pipeline_md_result[40]), .ZN(vscale_core_DW01_add_5n122) );
  NOR2_X2 vscale_core_DW01_add_5_U618 ( .A1(pipeline_md_b[43]), .A2(pipeline_md_result[43]), .ZN(vscale_core_DW01_add_5n105) );
  NOR2_X2 vscale_core_DW01_add_5_U619 ( .A1(pipeline_md_b[49]), .A2(pipeline_md_result[49]), .ZN(vscale_core_DW01_add_5n81) );
  NOR2_X2 vscale_core_DW01_add_5_U620 ( .A1(pipeline_md_b[47]), .A2(pipeline_md_result[47]), .ZN(vscale_core_DW01_add_5n89) );
  NOR2_X2 vscale_core_DW01_add_5_U621 ( .A1(pipeline_md_b[45]), .A2(pipeline_md_result[45]), .ZN(vscale_core_DW01_add_5n97) );
  OR2_X1 vscale_core_DW01_add_5_U622 ( .A1(pipeline_md_b[44]), .A2(pipeline_md_result[44]), .ZN(vscale_core_DW01_add_5n602) );
  OR2_X1 vscale_core_DW01_add_5_U623 ( .A1(pipeline_md_b[50]), .A2(pipeline_md_result[50]), .ZN(vscale_core_DW01_add_5n603) );
  OR2_X1 vscale_core_DW01_add_5_U624 ( .A1(pipeline_md_b[46]), .A2(pipeline_md_result[46]), .ZN(vscale_core_DW01_add_5n604) );
  OR2_X1 vscale_core_DW01_add_5_U625 ( .A1(pipeline_md_b[48]), .A2(pipeline_md_result[48]), .ZN(vscale_core_DW01_add_5n605) );
  NOR2_X2 vscale_core_DW01_add_5_U626 ( .A1(pipeline_md_b[53]), .A2(pipeline_md_result[53]), .ZN(vscale_core_DW01_add_5n65) );
  NOR2_X2 vscale_core_DW01_add_5_U627 ( .A1(pipeline_md_b[51]), .A2(pipeline_md_result[51]), .ZN(vscale_core_DW01_add_5n73) );
  OR2_X1 vscale_core_DW01_add_5_U628 ( .A1(pipeline_md_b[52]), .A2(pipeline_md_result[52]), .ZN(vscale_core_DW01_add_5n606) );
  OR2_X1 vscale_core_DW01_add_5_U629 ( .A1(pipeline_md_b[0]), .A2(pipeline_md_resp_result[0]), .ZN(vscale_core_DW01_add_5n607) );
  INV_X4 vscale_core_DW01_add_5_U630 ( .A(vscale_core_DW01_add_5n95), .ZN(vscale_core_DW01_add_5n93) );
  INV_X4 vscale_core_DW01_add_5_U631 ( .A(vscale_core_DW01_add_5n87), .ZN(vscale_core_DW01_add_5n85) );
  INV_X4 vscale_core_DW01_add_5_U632 ( .A(vscale_core_DW01_add_5n79), .ZN(vscale_core_DW01_add_5n77) );
  INV_X4 vscale_core_DW01_add_5_U633 ( .A(vscale_core_DW01_add_5n71), .ZN(vscale_core_DW01_add_5n69) );
  INV_X4 vscale_core_DW01_add_5_U634 ( .A(vscale_core_DW01_add_5n345), .ZN(vscale_core_DW01_add_5n401) );
  INV_X4 vscale_core_DW01_add_5_U635 ( .A(vscale_core_DW01_add_5n341), .ZN(vscale_core_DW01_add_5n400) );
  INV_X4 vscale_core_DW01_add_5_U636 ( .A(vscale_core_DW01_add_5n338), .ZN(vscale_core_DW01_add_5n399) );
  INV_X4 vscale_core_DW01_add_5_U637 ( .A(vscale_core_DW01_add_5n327), .ZN(vscale_core_DW01_add_5n397) );
  INV_X4 vscale_core_DW01_add_5_U638 ( .A(vscale_core_DW01_add_5n322), .ZN(vscale_core_DW01_add_5n396) );
  INV_X4 vscale_core_DW01_add_5_U639 ( .A(vscale_core_DW01_add_5n319), .ZN(vscale_core_DW01_add_5n395) );
  INV_X4 vscale_core_DW01_add_5_U640 ( .A(vscale_core_DW01_add_5n311), .ZN(vscale_core_DW01_add_5n394) );
  INV_X4 vscale_core_DW01_add_5_U641 ( .A(vscale_core_DW01_add_5n308), .ZN(vscale_core_DW01_add_5n393) );
  INV_X4 vscale_core_DW01_add_5_U642 ( .A(vscale_core_DW01_add_5n296), .ZN(vscale_core_DW01_add_5n391) );
  INV_X4 vscale_core_DW01_add_5_U643 ( .A(vscale_core_DW01_add_5n283), .ZN(vscale_core_DW01_add_5n389) );
  INV_X4 vscale_core_DW01_add_5_U644 ( .A(vscale_core_DW01_add_5n271), .ZN(vscale_core_DW01_add_5n387) );
  INV_X4 vscale_core_DW01_add_5_U645 ( .A(vscale_core_DW01_add_5n256), .ZN(vscale_core_DW01_add_5n385) );
  INV_X4 vscale_core_DW01_add_5_U646 ( .A(vscale_core_DW01_add_5n251), .ZN(vscale_core_DW01_add_5n384) );
  INV_X4 vscale_core_DW01_add_5_U647 ( .A(vscale_core_DW01_add_5n248), .ZN(vscale_core_DW01_add_5n383) );
  INV_X4 vscale_core_DW01_add_5_U648 ( .A(vscale_core_DW01_add_5n238), .ZN(vscale_core_DW01_add_5n382) );
  INV_X4 vscale_core_DW01_add_5_U649 ( .A(vscale_core_DW01_add_5n235), .ZN(vscale_core_DW01_add_5n381) );
  INV_X4 vscale_core_DW01_add_5_U650 ( .A(vscale_core_DW01_add_5n230), .ZN(vscale_core_DW01_add_5n380) );
  INV_X4 vscale_core_DW01_add_5_U651 ( .A(vscale_core_DW01_add_5n227), .ZN(vscale_core_DW01_add_5n379) );
  INV_X4 vscale_core_DW01_add_5_U652 ( .A(vscale_core_DW01_add_5n217), .ZN(vscale_core_DW01_add_5n378) );
  INV_X4 vscale_core_DW01_add_5_U653 ( .A(vscale_core_DW01_add_5n214), .ZN(vscale_core_DW01_add_5n377) );
  INV_X4 vscale_core_DW01_add_5_U654 ( .A(vscale_core_DW01_add_5n209), .ZN(vscale_core_DW01_add_5n376) );
  INV_X4 vscale_core_DW01_add_5_U655 ( .A(vscale_core_DW01_add_5n206), .ZN(vscale_core_DW01_add_5n375) );
  INV_X4 vscale_core_DW01_add_5_U656 ( .A(vscale_core_DW01_add_5n196), .ZN(vscale_core_DW01_add_5n374) );
  INV_X4 vscale_core_DW01_add_5_U657 ( .A(vscale_core_DW01_add_5n193), .ZN(vscale_core_DW01_add_5n373) );
  INV_X4 vscale_core_DW01_add_5_U658 ( .A(vscale_core_DW01_add_5n188), .ZN(vscale_core_DW01_add_5n372) );
  INV_X4 vscale_core_DW01_add_5_U659 ( .A(vscale_core_DW01_add_5n185), .ZN(vscale_core_DW01_add_5n371) );
  INV_X4 vscale_core_DW01_add_5_U660 ( .A(vscale_core_DW01_add_5n173), .ZN(vscale_core_DW01_add_5n370) );
  INV_X4 vscale_core_DW01_add_5_U661 ( .A(vscale_core_DW01_add_5n170), .ZN(vscale_core_DW01_add_5n369) );
  INV_X4 vscale_core_DW01_add_5_U662 ( .A(vscale_core_DW01_add_5n158), .ZN(vscale_core_DW01_add_5n367) );
  INV_X4 vscale_core_DW01_add_5_U663 ( .A(vscale_core_DW01_add_5n145), .ZN(vscale_core_DW01_add_5n365) );
  INV_X4 vscale_core_DW01_add_5_U664 ( .A(vscale_core_DW01_add_5n133), .ZN(vscale_core_DW01_add_5n363) );
  INV_X4 vscale_core_DW01_add_5_U665 ( .A(vscale_core_DW01_add_5n117), .ZN(vscale_core_DW01_add_5n361) );
  INV_X4 vscale_core_DW01_add_5_U666 ( .A(vscale_core_DW01_add_5n110), .ZN(vscale_core_DW01_add_5n360) );
  INV_X4 vscale_core_DW01_add_5_U667 ( .A(vscale_core_DW01_add_5n105), .ZN(vscale_core_DW01_add_5n359) );
  INV_X4 vscale_core_DW01_add_5_U668 ( .A(vscale_core_DW01_add_5n97), .ZN(vscale_core_DW01_add_5n357) );
  INV_X4 vscale_core_DW01_add_5_U669 ( .A(vscale_core_DW01_add_5n89), .ZN(vscale_core_DW01_add_5n355) );
  INV_X4 vscale_core_DW01_add_5_U670 ( .A(vscale_core_DW01_add_5n81), .ZN(vscale_core_DW01_add_5n353) );
  INV_X4 vscale_core_DW01_add_5_U671 ( .A(vscale_core_DW01_add_5n73), .ZN(vscale_core_DW01_add_5n351) );
  INV_X4 vscale_core_DW01_add_5_U672 ( .A(vscale_core_DW01_add_5n65), .ZN(vscale_core_DW01_add_5n349) );
  INV_X4 vscale_core_DW01_add_5_U673 ( .A(vscale_core_DW01_add_5n344), .ZN(vscale_core_DW01_add_5n343) );
  INV_X4 vscale_core_DW01_add_5_U674 ( .A(vscale_core_DW01_add_5n335), .ZN(vscale_core_DW01_add_5n334) );
  INV_X4 vscale_core_DW01_add_5_U675 ( .A(vscale_core_DW01_add_5n333), .ZN(vscale_core_DW01_add_5n331) );
  INV_X4 vscale_core_DW01_add_5_U676 ( .A(vscale_core_DW01_add_5n332), .ZN(vscale_core_DW01_add_5n398) );
  INV_X4 vscale_core_DW01_add_5_U677 ( .A(vscale_core_DW01_add_5n314), .ZN(vscale_core_DW01_add_5n313) );
  INV_X4 vscale_core_DW01_add_5_U678 ( .A(vscale_core_DW01_add_5n307), .ZN(vscale_core_DW01_add_5n305) );
  INV_X4 vscale_core_DW01_add_5_U679 ( .A(vscale_core_DW01_add_5n306), .ZN(vscale_core_DW01_add_5n304) );
  INV_X4 vscale_core_DW01_add_5_U680 ( .A(vscale_core_DW01_add_5n302), .ZN(vscale_core_DW01_add_5n300) );
  INV_X4 vscale_core_DW01_add_5_U681 ( .A(vscale_core_DW01_add_5n301), .ZN(vscale_core_DW01_add_5n392) );
  INV_X4 vscale_core_DW01_add_5_U682 ( .A(vscale_core_DW01_add_5n291), .ZN(vscale_core_DW01_add_5n290) );
  INV_X4 vscale_core_DW01_add_5_U683 ( .A(vscale_core_DW01_add_5n289), .ZN(vscale_core_DW01_add_5n287) );
  INV_X4 vscale_core_DW01_add_5_U684 ( .A(vscale_core_DW01_add_5n288), .ZN(vscale_core_DW01_add_5n390) );
  INV_X4 vscale_core_DW01_add_5_U685 ( .A(vscale_core_DW01_add_5n282), .ZN(vscale_core_DW01_add_5n280) );
  INV_X4 vscale_core_DW01_add_5_U686 ( .A(vscale_core_DW01_add_5n281), .ZN(vscale_core_DW01_add_5n279) );
  INV_X4 vscale_core_DW01_add_5_U687 ( .A(vscale_core_DW01_add_5n277), .ZN(vscale_core_DW01_add_5n275) );
  INV_X4 vscale_core_DW01_add_5_U688 ( .A(vscale_core_DW01_add_5n276), .ZN(vscale_core_DW01_add_5n388) );
  INV_X4 vscale_core_DW01_add_5_U689 ( .A(vscale_core_DW01_add_5n264), .ZN(vscale_core_DW01_add_5n263) );
  INV_X4 vscale_core_DW01_add_5_U690 ( .A(vscale_core_DW01_add_5n262), .ZN(vscale_core_DW01_add_5n260) );
  INV_X4 vscale_core_DW01_add_5_U691 ( .A(vscale_core_DW01_add_5n261), .ZN(vscale_core_DW01_add_5n386) );
  INV_X4 vscale_core_DW01_add_5_U692 ( .A(vscale_core_DW01_add_5n245), .ZN(vscale_core_DW01_add_5n243) );
  INV_X4 vscale_core_DW01_add_5_U693 ( .A(vscale_core_DW01_add_5n244), .ZN(vscale_core_DW01_add_5n242) );
  INV_X4 vscale_core_DW01_add_5_U694 ( .A(vscale_core_DW01_add_5n241), .ZN(vscale_core_DW01_add_5n240) );
  INV_X4 vscale_core_DW01_add_5_U695 ( .A(vscale_core_DW01_add_5n220), .ZN(vscale_core_DW01_add_5n219) );
  INV_X4 vscale_core_DW01_add_5_U696 ( .A(vscale_core_DW01_add_5n203), .ZN(vscale_core_DW01_add_5n201) );
  INV_X4 vscale_core_DW01_add_5_U697 ( .A(vscale_core_DW01_add_5n202), .ZN(vscale_core_DW01_add_5n200) );
  INV_X4 vscale_core_DW01_add_5_U698 ( .A(vscale_core_DW01_add_5n199), .ZN(vscale_core_DW01_add_5n198) );
  INV_X4 vscale_core_DW01_add_5_U699 ( .A(vscale_core_DW01_add_5n176), .ZN(vscale_core_DW01_add_5n175) );
  INV_X4 vscale_core_DW01_add_5_U700 ( .A(vscale_core_DW01_add_5n169), .ZN(vscale_core_DW01_add_5n167) );
  INV_X4 vscale_core_DW01_add_5_U701 ( .A(vscale_core_DW01_add_5n168), .ZN(vscale_core_DW01_add_5n166) );
  INV_X4 vscale_core_DW01_add_5_U702 ( .A(vscale_core_DW01_add_5n164), .ZN(vscale_core_DW01_add_5n162) );
  INV_X4 vscale_core_DW01_add_5_U703 ( .A(vscale_core_DW01_add_5n163), .ZN(vscale_core_DW01_add_5n368) );
  INV_X4 vscale_core_DW01_add_5_U704 ( .A(vscale_core_DW01_add_5n153), .ZN(vscale_core_DW01_add_5n152) );
  INV_X4 vscale_core_DW01_add_5_U705 ( .A(vscale_core_DW01_add_5n151), .ZN(vscale_core_DW01_add_5n149) );
  INV_X4 vscale_core_DW01_add_5_U706 ( .A(vscale_core_DW01_add_5n150), .ZN(vscale_core_DW01_add_5n366) );
  INV_X4 vscale_core_DW01_add_5_U707 ( .A(vscale_core_DW01_add_5n144), .ZN(vscale_core_DW01_add_5n142) );
  INV_X4 vscale_core_DW01_add_5_U708 ( .A(vscale_core_DW01_add_5n143), .ZN(vscale_core_DW01_add_5n141) );
  INV_X4 vscale_core_DW01_add_5_U709 ( .A(vscale_core_DW01_add_5n139), .ZN(vscale_core_DW01_add_5n137) );
  INV_X4 vscale_core_DW01_add_5_U710 ( .A(vscale_core_DW01_add_5n138), .ZN(vscale_core_DW01_add_5n364) );
  INV_X4 vscale_core_DW01_add_5_U711 ( .A(vscale_core_DW01_add_5n128), .ZN(vscale_core_DW01_add_5n126) );
  INV_X4 vscale_core_DW01_add_5_U712 ( .A(vscale_core_DW01_add_5n127), .ZN(vscale_core_DW01_add_5n125) );
  INV_X4 vscale_core_DW01_add_5_U713 ( .A(vscale_core_DW01_add_5n123), .ZN(vscale_core_DW01_add_5n121) );
  INV_X4 vscale_core_DW01_add_5_U714 ( .A(vscale_core_DW01_add_5n122), .ZN(vscale_core_DW01_add_5n362) );
  INV_X4 vscale_core_DW01_add_5_U715 ( .A(vscale_core_DW01_add_5n103), .ZN(vscale_core_DW01_add_5n101) );
;
  vscale_core_DW01_cmp6_1 r579 

  NAND2_X2 vscale_core_DW01_cmp6_1_U10 ( .A1(vscale_core_DW01_cmp6_1n36), .A2(vscale_core_DW01_cmp6_1n6), .ZN(vscale_core_DW01_cmp6_1n4) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U14 ( .A1(vscale_core_DW01_cmp6_1n16), .A2(vscale_core_DW01_cmp6_1n10), .ZN(vscale_core_DW01_cmp6_1n8) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U18 ( .A(vscale_core_DW01_cmp6_1n132), .B(pipeline_alu_N316), .ZN(vscale_core_DW01_cmp6_1n12) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U19 ( .A1(vscale_core_DW01_cmp6_1n132), .A2(pipeline_alu_N316), .ZN(vscale_core_DW01_cmp6_1n13) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U20 ( .A(vscale_core_DW01_cmp6_1n133), .B(pipeline_alu_src_a[30]), .ZN(vscale_core_DW01_cmp6_1n14) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U21 ( .A1(vscale_core_DW01_cmp6_1n133), .A2(pipeline_alu_src_a[30]), .ZN(vscale_core_DW01_cmp6_1n15) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U24 ( .A(vscale_core_DW01_cmp6_1n134), .B(pipeline_alu_src_a[29]), .ZN(vscale_core_DW01_cmp6_1n18) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U25 ( .A1(vscale_core_DW01_cmp6_1n134), .A2(pipeline_alu_src_a[29]), .ZN(vscale_core_DW01_cmp6_1n19) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U27 ( .A1(vscale_core_DW01_cmp6_1n135), .A2(n6563), .ZN(vscale_core_DW01_cmp6_1n21) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U32 ( .A(vscale_core_DW01_cmp6_1n136), .B(pipeline_alu_src_a[27]), .ZN(vscale_core_DW01_cmp6_1n26) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U34 ( .A(vscale_core_DW01_cmp6_1n137), .B(n6559), .ZN(vscale_core_DW01_cmp6_1n28) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U35 ( .A1(vscale_core_DW01_cmp6_1n137), .A2(n6559), .ZN(vscale_core_DW01_cmp6_1n29) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U38 ( .A(vscale_core_DW01_cmp6_1n138), .B(pipeline_alu_src_a[25]), .ZN(vscale_core_DW01_cmp6_1n32) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U40 ( .A(vscale_core_DW01_cmp6_1n139), .B(pipeline_alu_src_a[24]), .ZN(vscale_core_DW01_cmp6_1n34) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U41 ( .A1(vscale_core_DW01_cmp6_1n139), .A2(pipeline_alu_src_a[24]), .ZN(vscale_core_DW01_cmp6_1n35) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U44 ( .A1(vscale_core_DW01_cmp6_1n46), .A2(vscale_core_DW01_cmp6_1n40), .ZN(vscale_core_DW01_cmp6_1n38) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U48 ( .A(vscale_core_DW01_cmp6_1n140), .B(pipeline_alu_src_a[23]), .ZN(vscale_core_DW01_cmp6_1n42) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U50 ( .A(vscale_core_DW01_cmp6_1n141), .B(pipeline_alu_src_a[22]), .ZN(vscale_core_DW01_cmp6_1n44) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U54 ( .A(vscale_core_DW01_cmp6_1n142), .B(pipeline_alu_src_a[21]), .ZN(vscale_core_DW01_cmp6_1n48) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U55 ( .A1(vscale_core_DW01_cmp6_1n142), .A2(pipeline_alu_src_a[21]), .ZN(vscale_core_DW01_cmp6_1n49) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U57 ( .A1(vscale_core_DW01_cmp6_1n143), .A2(pipeline_alu_src_a[20]), .ZN(vscale_core_DW01_cmp6_1n51) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U58 ( .A1(vscale_core_DW01_cmp6_1n60), .A2(vscale_core_DW01_cmp6_1n54), .ZN(vscale_core_DW01_cmp6_1n52) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U63 ( .A1(vscale_core_DW01_cmp6_1n144), .A2(pipeline_alu_src_a[19]), .ZN(vscale_core_DW01_cmp6_1n57) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U64 ( .A(vscale_core_DW01_cmp6_1n145), .B(pipeline_alu_src_a[18]), .ZN(vscale_core_DW01_cmp6_1n58) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U68 ( .A(vscale_core_DW01_cmp6_1n146), .B(pipeline_alu_src_a[17]), .ZN(vscale_core_DW01_cmp6_1n62) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U82 ( .A(vscale_core_DW01_cmp6_1n149), .B(pipeline_alu_src_a[14]), .ZN(vscale_core_DW01_cmp6_1n76) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U83 ( .A1(vscale_core_DW01_cmp6_1n149), .A2(pipeline_alu_src_a[14]), .ZN(vscale_core_DW01_cmp6_1n77) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U86 ( .A(vscale_core_DW01_cmp6_1n150), .B(n6568), .ZN(vscale_core_DW01_cmp6_1n80) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U87 ( .A1(vscale_core_DW01_cmp6_1n150), .A2(n6568), .ZN(vscale_core_DW01_cmp6_1n81) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U90 ( .A1(vscale_core_DW01_cmp6_1n92), .A2(vscale_core_DW01_cmp6_1n86), .ZN(vscale_core_DW01_cmp6_1n84) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U100 ( .A(vscale_core_DW01_cmp6_1n154), .B(n6973), .ZN(vscale_core_DW01_cmp6_1n94) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U101 ( .A1(vscale_core_DW01_cmp6_1n154), .A2(n6973), .ZN(vscale_core_DW01_cmp6_1n95) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U106 ( .A1(vscale_core_DW01_cmp6_1n108), .A2(vscale_core_DW01_cmp6_1n102), .ZN(vscale_core_DW01_cmp6_1n100) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U120 ( .A1(vscale_core_DW01_cmp6_1n116), .A2(vscale_core_DW01_cmp6_1n122), .ZN(vscale_core_DW01_cmp6_1n114) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U124 ( .A(vscale_core_DW01_cmp6_1n160), .B(n6635), .ZN(vscale_core_DW01_cmp6_1n118) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U130 ( .A(vscale_core_DW01_cmp6_1n162), .B(n6632), .ZN(vscale_core_DW01_cmp6_1n124) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U131 ( .A1(vscale_core_DW01_cmp6_1n162), .A2(n6632), .ZN(vscale_core_DW01_cmp6_1n125) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U173 ( .A1(vscale_core_DW01_cmp6_1n28), .A2(vscale_core_DW01_cmp6_1n26), .ZN(vscale_core_DW01_cmp6_1n24) );
  INV_X2 vscale_core_DW01_cmp6_1_U174 ( .A(pipeline_alu_src_b[8]), .ZN(vscale_core_DW01_cmp6_1n155) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U175 ( .A1(vscale_core_DW01_cmp6_1n22), .A2(vscale_core_DW01_cmp6_1n8), .ZN(vscale_core_DW01_cmp6_1n6) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U176 ( .B1(vscale_core_DW01_cmp6_1n37), .B2(vscale_core_DW01_cmp6_1n6), .A(vscale_core_DW01_cmp6_1n7), .ZN(vscale_core_DW01_cmp6_1n5) );
  INV_X1 vscale_core_DW01_cmp6_1_U177 ( .A(pipeline_alu_src_b[7]), .ZN(vscale_core_DW01_cmp6_1n156) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U178 ( .A1(vscale_core_DW01_cmp6_1n76), .A2(vscale_core_DW01_cmp6_1n74), .ZN(vscale_core_DW01_cmp6_1n72) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U179 ( .A1(vscale_core_DW01_cmp6_1n104), .A2(vscale_core_DW01_cmp6_1n106), .ZN(vscale_core_DW01_cmp6_1n102) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U180 ( .B1(vscale_core_DW01_cmp6_1n118), .B2(vscale_core_DW01_cmp6_1n121), .A(vscale_core_DW01_cmp6_1n119), .ZN(vscale_core_DW01_cmp6_1n117) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U181 ( .B1(vscale_core_DW01_cmp6_1n54), .B2(vscale_core_DW01_cmp6_1n61), .A(vscale_core_DW01_cmp6_1n55), .ZN(vscale_core_DW01_cmp6_1n53) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U182 ( .B1(vscale_core_DW01_cmp6_1n56), .B2(vscale_core_DW01_cmp6_1n59), .A(vscale_core_DW01_cmp6_1n57), .ZN(vscale_core_DW01_cmp6_1n55) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U183 ( .B1(vscale_core_DW01_cmp6_1n102), .B2(vscale_core_DW01_cmp6_1n109), .A(vscale_core_DW01_cmp6_1n103), .ZN(vscale_core_DW01_cmp6_1n101) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U184 ( .B1(vscale_core_DW01_cmp6_1n110), .B2(vscale_core_DW01_cmp6_1n113), .A(vscale_core_DW01_cmp6_1n111), .ZN(vscale_core_DW01_cmp6_1n109) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U185 ( .B1(vscale_core_DW01_cmp6_1n72), .B2(vscale_core_DW01_cmp6_1n79), .A(vscale_core_DW01_cmp6_1n73), .ZN(vscale_core_DW01_cmp6_1n71) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U186 ( .A1(vscale_core_DW01_cmp6_1n120), .A2(vscale_core_DW01_cmp6_1n118), .ZN(vscale_core_DW01_cmp6_1n116) );
  NOR2_X1 vscale_core_DW01_cmp6_1_U187 ( .A1(vscale_core_DW01_cmp6_1n52), .A2(vscale_core_DW01_cmp6_1n38), .ZN(vscale_core_DW01_cmp6_1n36) );
  NOR2_X1 vscale_core_DW01_cmp6_1_U188 ( .A1(vscale_core_DW01_cmp6_1n64), .A2(vscale_core_DW01_cmp6_1n62), .ZN(vscale_core_DW01_cmp6_1n60) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U189 ( .A1(vscale_core_DW01_cmp6_1n128), .A2(vscale_core_DW01_cmp6_1n240), .ZN(vscale_core_DW01_cmp6_1n127) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U190 ( .A1(vscale_core_DW01_cmp6_1n44), .A2(vscale_core_DW01_cmp6_1n42), .ZN(vscale_core_DW01_cmp6_1n40) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U191 ( .B1(vscale_core_DW01_cmp6_1n32), .B2(vscale_core_DW01_cmp6_1n35), .A(vscale_core_DW01_cmp6_1n33), .ZN(vscale_core_DW01_cmp6_1n31) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U192 ( .B1(vscale_core_DW01_cmp6_1n17), .B2(vscale_core_DW01_cmp6_1n10), .A(vscale_core_DW01_cmp6_1n11), .ZN(vscale_core_DW01_cmp6_1n9) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U193 ( .B1(vscale_core_DW01_cmp6_1n18), .B2(vscale_core_DW01_cmp6_1n21), .A(vscale_core_DW01_cmp6_1n19), .ZN(vscale_core_DW01_cmp6_1n17) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U194 ( .A1(vscale_core_DW01_cmp6_1n58), .A2(vscale_core_DW01_cmp6_1n56), .ZN(vscale_core_DW01_cmp6_1n54) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U195 ( .B1(vscale_core_DW01_cmp6_1n99), .B2(vscale_core_DW01_cmp6_1n68), .A(vscale_core_DW01_cmp6_1n69), .ZN(vscale_core_DW01_cmp6_1n67) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U196 ( .B1(vscale_core_DW01_cmp6_1n86), .B2(vscale_core_DW01_cmp6_1n93), .A(vscale_core_DW01_cmp6_1n87), .ZN(vscale_core_DW01_cmp6_1n85) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U197 ( .A1(vscale_core_DW01_cmp6_1n4), .A2(vscale_core_DW01_cmp6_1n66), .ZN(pipeline_alu_N251) );
  AND2_X4 vscale_core_DW01_cmp6_1_U198 ( .A1(vscale_core_DW01_cmp6_1n163), .A2(pipeline_alu_src_a[0]), .ZN(vscale_core_DW01_cmp6_1n240) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U199 ( .B1(vscale_core_DW01_cmp6_1n80), .B2(vscale_core_DW01_cmp6_1n83), .A(vscale_core_DW01_cmp6_1n81), .ZN(vscale_core_DW01_cmp6_1n79) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U200 ( .B1(vscale_core_DW01_cmp6_1n48), .B2(vscale_core_DW01_cmp6_1n51), .A(vscale_core_DW01_cmp6_1n49), .ZN(vscale_core_DW01_cmp6_1n47) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U201 ( .A1(vscale_core_DW01_cmp6_1n136), .A2(pipeline_alu_src_a[27]), .ZN(vscale_core_DW01_cmp6_1n27) );
  INV_X2 vscale_core_DW01_cmp6_1_U202 ( .A(pipeline_alu_src_b[15]), .ZN(vscale_core_DW01_cmp6_1n148) );
  INV_X1 vscale_core_DW01_cmp6_1_U203 ( .A(pipeline_alu_src_b[12]), .ZN(vscale_core_DW01_cmp6_1n151) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U204 ( .A1(vscale_core_DW01_cmp6_1n144), .A2(pipeline_alu_src_a[19]), .ZN(vscale_core_DW01_cmp6_1n242) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U205 ( .A1(pipeline_alu_src_b[19]), .A2(vscale_core_DW01_cmp6_1n241), .ZN(vscale_core_DW01_cmp6_1n243) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U206 ( .A1(vscale_core_DW01_cmp6_1n242), .A2(vscale_core_DW01_cmp6_1n243), .ZN(vscale_core_DW01_cmp6_1n56) );
  INV_X4 vscale_core_DW01_cmp6_1_U207 ( .A(pipeline_alu_src_a[19]), .ZN(vscale_core_DW01_cmp6_1n241) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U208 ( .A1(vscale_core_DW01_cmp6_1n140), .A2(pipeline_alu_src_a[23]), .ZN(vscale_core_DW01_cmp6_1n43) );
  INV_X2 vscale_core_DW01_cmp6_1_U209 ( .A(pipeline_alu_src_b[16]), .ZN(vscale_core_DW01_cmp6_1n147) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U210 ( .B1(vscale_core_DW01_cmp6_1n23), .B2(vscale_core_DW01_cmp6_1n8), .A(vscale_core_DW01_cmp6_1n9), .ZN(vscale_core_DW01_cmp6_1n7) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U211 ( .B1(vscale_core_DW01_cmp6_1n24), .B2(vscale_core_DW01_cmp6_1n31), .A(vscale_core_DW01_cmp6_1n25), .ZN(vscale_core_DW01_cmp6_1n23) );
  OAI21_X1 vscale_core_DW01_cmp6_1_U212 ( .B1(vscale_core_DW01_cmp6_1n12), .B2(vscale_core_DW01_cmp6_1n15), .A(vscale_core_DW01_cmp6_1n13), .ZN(vscale_core_DW01_cmp6_1n11) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U213 ( .A1(vscale_core_DW01_cmp6_1n156), .A2(n6612), .ZN(vscale_core_DW01_cmp6_1n105) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U214 ( .A(vscale_core_DW01_cmp6_1n156), .B(n6612), .ZN(vscale_core_DW01_cmp6_1n104) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U215 ( .A1(vscale_core_DW01_cmp6_1n30), .A2(vscale_core_DW01_cmp6_1n24), .ZN(vscale_core_DW01_cmp6_1n22) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U216 ( .A1(vscale_core_DW01_cmp6_1n14), .A2(vscale_core_DW01_cmp6_1n12), .ZN(vscale_core_DW01_cmp6_1n10) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U217 ( .A(vscale_core_DW01_cmp6_1n158), .B(n6620), .ZN(vscale_core_DW01_cmp6_1n110) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U218 ( .A1(vscale_core_DW01_cmp6_1n161), .A2(pipeline_alu_src_a[2]), .ZN(vscale_core_DW01_cmp6_1n121) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U219 ( .A(vscale_core_DW01_cmp6_1n161), .B(pipeline_alu_src_a[2]), .ZN(vscale_core_DW01_cmp6_1n120) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U220 ( .A(vscale_core_DW01_cmp6_1n163), .B(pipeline_alu_src_a[0]), .ZN(vscale_core_DW01_cmp6_1n126) );
  INV_X2 vscale_core_DW01_cmp6_1_U221 ( .A(pipeline_alu_src_b[5]), .ZN(vscale_core_DW01_cmp6_1n158) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U222 ( .A1(vscale_core_DW01_cmp6_1n152), .A2(pipeline_alu_src_a[11]), .ZN(vscale_core_DW01_cmp6_1n89) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U223 ( .A(vscale_core_DW01_cmp6_1n152), .B(pipeline_alu_src_a[11]), .ZN(vscale_core_DW01_cmp6_1n88) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U224 ( .A1(vscale_core_DW01_cmp6_1n146), .A2(pipeline_alu_src_a[17]), .ZN(vscale_core_DW01_cmp6_1n63) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U225 ( .A1(vscale_core_DW01_cmp6_1n98), .A2(vscale_core_DW01_cmp6_1n68), .ZN(vscale_core_DW01_cmp6_1n66) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U226 ( .A1(vscale_core_DW01_cmp6_1n70), .A2(vscale_core_DW01_cmp6_1n84), .ZN(vscale_core_DW01_cmp6_1n68) );
  NOR2_X1 vscale_core_DW01_cmp6_1_U227 ( .A1(vscale_core_DW01_cmp6_1n94), .A2(vscale_core_DW01_cmp6_1n96), .ZN(vscale_core_DW01_cmp6_1n92) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U228 ( .A1(vscale_core_DW01_cmp6_1n158), .A2(n6620), .ZN(vscale_core_DW01_cmp6_1n111) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U229 ( .A1(vscale_core_DW01_cmp6_1n159), .A2(n6928), .ZN(vscale_core_DW01_cmp6_1n113) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U230 ( .B1(vscale_core_DW01_cmp6_1n26), .B2(vscale_core_DW01_cmp6_1n29), .A(vscale_core_DW01_cmp6_1n27), .ZN(vscale_core_DW01_cmp6_1n25) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U231 ( .A1(vscale_core_DW01_cmp6_1n112), .A2(vscale_core_DW01_cmp6_1n110), .ZN(vscale_core_DW01_cmp6_1n108) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U232 ( .A(vscale_core_DW01_cmp6_1n135), .B(n6563), .ZN(vscale_core_DW01_cmp6_1n20) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U233 ( .B1(vscale_core_DW01_cmp6_1n42), .B2(vscale_core_DW01_cmp6_1n45), .A(vscale_core_DW01_cmp6_1n43), .ZN(vscale_core_DW01_cmp6_1n41) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U234 ( .A1(vscale_core_DW01_cmp6_1n141), .A2(pipeline_alu_src_a[22]), .ZN(vscale_core_DW01_cmp6_1n45) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U235 ( .A1(vscale_core_DW01_cmp6_1n138), .A2(pipeline_alu_src_a[25]), .ZN(vscale_core_DW01_cmp6_1n33) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U236 ( .A1(vscale_core_DW01_cmp6_1n145), .A2(pipeline_alu_src_a[18]), .ZN(vscale_core_DW01_cmp6_1n59) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U237 ( .A(vscale_core_DW01_cmp6_1n143), .B(pipeline_alu_src_a[20]), .ZN(vscale_core_DW01_cmp6_1n50) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U238 ( .A(vscale_core_DW01_cmp6_1n159), .B(n6928), .ZN(vscale_core_DW01_cmp6_1n112) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U239 ( .B1(vscale_core_DW01_cmp6_1n123), .B2(vscale_core_DW01_cmp6_1n116), .A(vscale_core_DW01_cmp6_1n117), .ZN(vscale_core_DW01_cmp6_1n115) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U240 ( .B1(vscale_core_DW01_cmp6_1n104), .B2(vscale_core_DW01_cmp6_1n107), .A(vscale_core_DW01_cmp6_1n105), .ZN(vscale_core_DW01_cmp6_1n103) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U241 ( .B1(vscale_core_DW01_cmp6_1n94), .B2(vscale_core_DW01_cmp6_1n97), .A(vscale_core_DW01_cmp6_1n95), .ZN(vscale_core_DW01_cmp6_1n93) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U242 ( .B1(vscale_core_DW01_cmp6_1n53), .B2(vscale_core_DW01_cmp6_1n38), .A(vscale_core_DW01_cmp6_1n39), .ZN(vscale_core_DW01_cmp6_1n37) );
  AOI21_X2 vscale_core_DW01_cmp6_1_U243 ( .B1(vscale_core_DW01_cmp6_1n40), .B2(vscale_core_DW01_cmp6_1n47), .A(vscale_core_DW01_cmp6_1n41), .ZN(vscale_core_DW01_cmp6_1n39) );
  NOR2_X1 vscale_core_DW01_cmp6_1_U244 ( .A1(vscale_core_DW01_cmp6_1n114), .A2(vscale_core_DW01_cmp6_1n100), .ZN(vscale_core_DW01_cmp6_1n98) );
  NOR2_X1 vscale_core_DW01_cmp6_1_U245 ( .A1(vscale_core_DW01_cmp6_1n126), .A2(vscale_core_DW01_cmp6_1n124), .ZN(vscale_core_DW01_cmp6_1n122) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U246 ( .B1(vscale_core_DW01_cmp6_1n62), .B2(vscale_core_DW01_cmp6_1n65), .A(vscale_core_DW01_cmp6_1n63), .ZN(vscale_core_DW01_cmp6_1n61) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U247 ( .A1(vscale_core_DW01_cmp6_1n50), .A2(vscale_core_DW01_cmp6_1n48), .ZN(vscale_core_DW01_cmp6_1n46) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U248 ( .B1(vscale_core_DW01_cmp6_1n127), .B2(vscale_core_DW01_cmp6_1n124), .A(vscale_core_DW01_cmp6_1n125), .ZN(vscale_core_DW01_cmp6_1n123) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U249 ( .B1(vscale_core_DW01_cmp6_1n88), .B2(vscale_core_DW01_cmp6_1n91), .A(vscale_core_DW01_cmp6_1n89), .ZN(vscale_core_DW01_cmp6_1n87) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U250 ( .A1(vscale_core_DW01_cmp6_1n20), .A2(vscale_core_DW01_cmp6_1n18), .ZN(vscale_core_DW01_cmp6_1n16) );
  NOR2_X1 vscale_core_DW01_cmp6_1_U251 ( .A1(vscale_core_DW01_cmp6_1n88), .A2(vscale_core_DW01_cmp6_1n90), .ZN(vscale_core_DW01_cmp6_1n86) );
  NOR2_X1 vscale_core_DW01_cmp6_1_U252 ( .A1(vscale_core_DW01_cmp6_1n34), .A2(vscale_core_DW01_cmp6_1n32), .ZN(vscale_core_DW01_cmp6_1n30) );
  NAND2_X2 vscale_core_DW01_cmp6_1_U253 ( .A1(vscale_core_DW01_cmp6_1n78), .A2(vscale_core_DW01_cmp6_1n72), .ZN(vscale_core_DW01_cmp6_1n70) );
  NOR2_X2 vscale_core_DW01_cmp6_1_U254 ( .A1(vscale_core_DW01_cmp6_1n82), .A2(vscale_core_DW01_cmp6_1n80), .ZN(vscale_core_DW01_cmp6_1n78) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U255 ( .A1(vscale_core_DW01_cmp6_1n153), .A2(n6572), .ZN(vscale_core_DW01_cmp6_1n91) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U256 ( .A(vscale_core_DW01_cmp6_1n153), .B(n6572), .ZN(vscale_core_DW01_cmp6_1n90) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U257 ( .A1(vscale_core_DW01_cmp6_1n151), .A2(pipeline_alu_src_a[12]), .ZN(vscale_core_DW01_cmp6_1n83) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U258 ( .A(vscale_core_DW01_cmp6_1n151), .B(pipeline_alu_src_a[12]), .ZN(vscale_core_DW01_cmp6_1n82) );
  INV_X2 vscale_core_DW01_cmp6_1_U259 ( .A(n6976), .ZN(vscale_core_DW01_cmp6_1n162) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U260 ( .A1(vscale_core_DW01_cmp6_1n148), .A2(n6598), .ZN(vscale_core_DW01_cmp6_1n75) );
  XNOR2_X2 vscale_core_DW01_cmp6_1_U261 ( .A(vscale_core_DW01_cmp6_1n148), .B(n6598), .ZN(vscale_core_DW01_cmp6_1n74) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U262 ( .A(vscale_core_DW01_cmp6_1n147), .B(pipeline_alu_src_a[16]), .ZN(vscale_core_DW01_cmp6_1n64) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U263 ( .A1(vscale_core_DW01_cmp6_1n147), .A2(pipeline_alu_src_a[16]), .ZN(vscale_core_DW01_cmp6_1n65) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U264 ( .A1(vscale_core_DW01_cmp6_1n157), .A2(n6605), .ZN(vscale_core_DW01_cmp6_1n107) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U265 ( .A(vscale_core_DW01_cmp6_1n157), .B(n6605), .ZN(vscale_core_DW01_cmp6_1n106) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U266 ( .B1(vscale_core_DW01_cmp6_1n74), .B2(vscale_core_DW01_cmp6_1n77), .A(vscale_core_DW01_cmp6_1n75), .ZN(vscale_core_DW01_cmp6_1n73) );
  OAI21_X4 vscale_core_DW01_cmp6_1_U267 ( .B1(vscale_core_DW01_cmp6_1n67), .B2(vscale_core_DW01_cmp6_1n4), .A(vscale_core_DW01_cmp6_1n5), .ZN(        pipeline_alu_N320) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U268 ( .A1(vscale_core_DW01_cmp6_1n155), .A2(n9335), .ZN(vscale_core_DW01_cmp6_1n97) );
  XNOR2_X1 vscale_core_DW01_cmp6_1_U269 ( .A(vscale_core_DW01_cmp6_1n155), .B(n9335), .ZN(vscale_core_DW01_cmp6_1n96) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U270 ( .B1(vscale_core_DW01_cmp6_1n85), .B2(vscale_core_DW01_cmp6_1n70), .A(vscale_core_DW01_cmp6_1n71), .ZN(vscale_core_DW01_cmp6_1n69) );
  OAI21_X2 vscale_core_DW01_cmp6_1_U271 ( .B1(vscale_core_DW01_cmp6_1n115), .B2(vscale_core_DW01_cmp6_1n100), .A(vscale_core_DW01_cmp6_1n101), .ZN(vscale_core_DW01_cmp6_1n99) );
  NAND2_X1 vscale_core_DW01_cmp6_1_U272 ( .A1(vscale_core_DW01_cmp6_1n160), .A2(n6635), .ZN(vscale_core_DW01_cmp6_1n119) );
  INV_X2 vscale_core_DW01_cmp6_1_U273 ( .A(n9339), .ZN(vscale_core_DW01_cmp6_1n160) );
  INV_X4 vscale_core_DW01_cmp6_1_U274 ( .A(n6618), .ZN(vscale_core_DW01_cmp6_1n163) );
  INV_X4 vscale_core_DW01_cmp6_1_U275 ( .A(n9398), .ZN(vscale_core_DW01_cmp6_1n161) );
  INV_X4 vscale_core_DW01_cmp6_1_U276 ( .A(pipeline_alu_src_b[4]), .ZN(vscale_core_DW01_cmp6_1n159) );
  INV_X4 vscale_core_DW01_cmp6_1_U277 ( .A(pipeline_alu_src_b[6]), .ZN(vscale_core_DW01_cmp6_1n157) );
  INV_X4 vscale_core_DW01_cmp6_1_U278 ( .A(pipeline_alu_src_b[9]), .ZN(vscale_core_DW01_cmp6_1n154) );
  INV_X4 vscale_core_DW01_cmp6_1_U279 ( .A(pipeline_alu_src_b[10]), .ZN(vscale_core_DW01_cmp6_1n153) );
  INV_X4 vscale_core_DW01_cmp6_1_U280 ( .A(pipeline_alu_src_b[11]), .ZN(vscale_core_DW01_cmp6_1n152) );
  INV_X4 vscale_core_DW01_cmp6_1_U281 ( .A(pipeline_alu_src_b[13]), .ZN(vscale_core_DW01_cmp6_1n150) );
  INV_X4 vscale_core_DW01_cmp6_1_U282 ( .A(pipeline_alu_src_b[14]), .ZN(vscale_core_DW01_cmp6_1n149) );
  INV_X4 vscale_core_DW01_cmp6_1_U283 ( .A(pipeline_alu_src_b[17]), .ZN(vscale_core_DW01_cmp6_1n146) );
  INV_X4 vscale_core_DW01_cmp6_1_U284 ( .A(pipeline_alu_src_b[18]), .ZN(vscale_core_DW01_cmp6_1n145) );
  INV_X4 vscale_core_DW01_cmp6_1_U285 ( .A(pipeline_alu_src_b[19]), .ZN(vscale_core_DW01_cmp6_1n144) );
  INV_X4 vscale_core_DW01_cmp6_1_U286 ( .A(pipeline_alu_src_b[20]), .ZN(vscale_core_DW01_cmp6_1n143) );
  INV_X4 vscale_core_DW01_cmp6_1_U287 ( .A(pipeline_alu_src_b[21]), .ZN(vscale_core_DW01_cmp6_1n142) );
  INV_X4 vscale_core_DW01_cmp6_1_U288 ( .A(pipeline_alu_src_b[22]), .ZN(vscale_core_DW01_cmp6_1n141) );
  INV_X4 vscale_core_DW01_cmp6_1_U289 ( .A(pipeline_alu_src_b[23]), .ZN(vscale_core_DW01_cmp6_1n140) );
  INV_X4 vscale_core_DW01_cmp6_1_U290 ( .A(pipeline_alu_src_b[24]), .ZN(vscale_core_DW01_cmp6_1n139) );
  INV_X4 vscale_core_DW01_cmp6_1_U291 ( .A(pipeline_alu_src_b[25]), .ZN(vscale_core_DW01_cmp6_1n138) );
  INV_X4 vscale_core_DW01_cmp6_1_U292 ( .A(pipeline_alu_src_b[26]), .ZN(vscale_core_DW01_cmp6_1n137) );
  INV_X4 vscale_core_DW01_cmp6_1_U293 ( .A(pipeline_alu_src_b[27]), .ZN(vscale_core_DW01_cmp6_1n136) );
  INV_X4 vscale_core_DW01_cmp6_1_U294 ( .A(pipeline_alu_src_b[28]), .ZN(vscale_core_DW01_cmp6_1n135) );
  INV_X4 vscale_core_DW01_cmp6_1_U295 ( .A(pipeline_alu_src_b[29]), .ZN(vscale_core_DW01_cmp6_1n134) );
  INV_X4 vscale_core_DW01_cmp6_1_U296 ( .A(pipeline_alu_src_b[30]), .ZN(vscale_core_DW01_cmp6_1n133) );
  INV_X4 vscale_core_DW01_cmp6_1_U297 ( .A(n13159), .ZN(vscale_core_DW01_cmp6_1n132) );
  INV_X4 vscale_core_DW01_cmp6_1_U298 ( .A(vscale_core_DW01_cmp6_1n126), .ZN(vscale_core_DW01_cmp6_1n128) );
  INV_X4 vscale_core_DW01_cmp6_1_U299 ( .A(pipeline_alu_N251), .ZN(pipeline_alu_N252) );
  INV_X4 vscale_core_DW01_cmp6_1_U300 ( .A(        pipeline_alu_N320), .ZN(pipeline_alu_N319) );
;
  vscale_core_DW01_sub_7 pipeline_alu_sub_25 

  XOR2_X2 vscale_core_DW01_sub_7_U1 ( .A(vscale_core_DW01_sub_7n1), .B(vscale_core_DW01_sub_7n29), .Z(pipeline_alu_N284) );
  FA_X1 vscale_core_DW01_sub_7_U3 ( .A(vscale_core_DW01_sub_7n206), .B(n6997), .CI(vscale_core_DW01_sub_7n30), .CO(vscale_core_DW01_sub_7n29), .S(pipeline_alu_N283) );
  FA_X1 vscale_core_DW01_sub_7_U4 ( .A(vscale_core_DW01_sub_7n207), .B(pipeline_alu_src_a[29]), .CI(vscale_core_DW01_sub_7n31), .CO(vscale_core_DW01_sub_7n30), .S(pipeline_alu_N282) );
  FA_X1 vscale_core_DW01_sub_7_U5 ( .A(vscale_core_DW01_sub_7n208), .B(n6564), .CI(vscale_core_DW01_sub_7n177), .CO(vscale_core_DW01_sub_7n31), .S(pipeline_alu_N281) );
  XNOR2_X2 vscale_core_DW01_sub_7_U7 ( .A(vscale_core_DW01_sub_7n37), .B(vscale_core_DW01_sub_7n2), .ZN(pipeline_alu_N280) );
  NAND2_X2 vscale_core_DW01_sub_7_U11 ( .A1(vscale_core_DW01_sub_7n343), .A2(vscale_core_DW01_sub_7n36), .ZN(vscale_core_DW01_sub_7n2) );
  XOR2_X2 vscale_core_DW01_sub_7_U15 ( .A(vscale_core_DW01_sub_7n3), .B(vscale_core_DW01_sub_7n40), .Z(pipeline_alu_N279) );
  NAND2_X2 vscale_core_DW01_sub_7_U17 ( .A1(vscale_core_DW01_sub_7n179), .A2(vscale_core_DW01_sub_7n39), .ZN(vscale_core_DW01_sub_7n3) );
  NAND2_X2 vscale_core_DW01_sub_7_U20 ( .A1(vscale_core_DW01_sub_7n210), .A2(n6561), .ZN(vscale_core_DW01_sub_7n39) );
  XNOR2_X2 vscale_core_DW01_sub_7_U21 ( .A(vscale_core_DW01_sub_7n45), .B(vscale_core_DW01_sub_7n4), .ZN(pipeline_alu_N278) );
  NAND2_X2 vscale_core_DW01_sub_7_U25 ( .A1(vscale_core_DW01_sub_7n344), .A2(vscale_core_DW01_sub_7n44), .ZN(vscale_core_DW01_sub_7n4) );
  NAND2_X2 vscale_core_DW01_sub_7_U28 ( .A1(vscale_core_DW01_sub_7n211), .A2(n6609), .ZN(vscale_core_DW01_sub_7n44) );
  XOR2_X2 vscale_core_DW01_sub_7_U29 ( .A(vscale_core_DW01_sub_7n5), .B(vscale_core_DW01_sub_7n48), .Z(pipeline_alu_N277) );
  NAND2_X2 vscale_core_DW01_sub_7_U31 ( .A1(vscale_core_DW01_sub_7n181), .A2(vscale_core_DW01_sub_7n47), .ZN(vscale_core_DW01_sub_7n5) );
  NAND2_X2 vscale_core_DW01_sub_7_U34 ( .A1(vscale_core_DW01_sub_7n212), .A2(pipeline_alu_src_a[24]), .ZN(vscale_core_DW01_sub_7n47) );
  XNOR2_X2 vscale_core_DW01_sub_7_U35 ( .A(vscale_core_DW01_sub_7n53), .B(vscale_core_DW01_sub_7n6), .ZN(pipeline_alu_N276) );
  NAND2_X2 vscale_core_DW01_sub_7_U39 ( .A1(vscale_core_DW01_sub_7n342), .A2(vscale_core_DW01_sub_7n52), .ZN(vscale_core_DW01_sub_7n6) );
  NAND2_X2 vscale_core_DW01_sub_7_U42 ( .A1(vscale_core_DW01_sub_7n213), .A2(n6980), .ZN(vscale_core_DW01_sub_7n52) );
  XOR2_X2 vscale_core_DW01_sub_7_U43 ( .A(vscale_core_DW01_sub_7n7), .B(vscale_core_DW01_sub_7n56), .Z(pipeline_alu_N275) );
  NAND2_X2 vscale_core_DW01_sub_7_U45 ( .A1(vscale_core_DW01_sub_7n183), .A2(vscale_core_DW01_sub_7n55), .ZN(vscale_core_DW01_sub_7n7) );
  NAND2_X2 vscale_core_DW01_sub_7_U48 ( .A1(vscale_core_DW01_sub_7n214), .A2(n6625), .ZN(vscale_core_DW01_sub_7n55) );
  XNOR2_X2 vscale_core_DW01_sub_7_U49 ( .A(vscale_core_DW01_sub_7n61), .B(vscale_core_DW01_sub_7n8), .ZN(pipeline_alu_N274) );
  NAND2_X2 vscale_core_DW01_sub_7_U53 ( .A1(vscale_core_DW01_sub_7n341), .A2(vscale_core_DW01_sub_7n60), .ZN(vscale_core_DW01_sub_7n8) );
  NAND2_X2 vscale_core_DW01_sub_7_U56 ( .A1(vscale_core_DW01_sub_7n215), .A2(pipeline_alu_src_a[21]), .ZN(vscale_core_DW01_sub_7n60) );
  XOR2_X2 vscale_core_DW01_sub_7_U57 ( .A(vscale_core_DW01_sub_7n9), .B(vscale_core_DW01_sub_7n68), .Z(pipeline_alu_N273) );
  NAND2_X2 vscale_core_DW01_sub_7_U59 ( .A1(vscale_core_DW01_sub_7n69), .A2(vscale_core_DW01_sub_7n340), .ZN(vscale_core_DW01_sub_7n62) );
  NAND2_X2 vscale_core_DW01_sub_7_U63 ( .A1(vscale_core_DW01_sub_7n340), .A2(vscale_core_DW01_sub_7n67), .ZN(vscale_core_DW01_sub_7n9) );
  NAND2_X2 vscale_core_DW01_sub_7_U66 ( .A1(vscale_core_DW01_sub_7n216), .A2(pipeline_alu_src_a[20]), .ZN(vscale_core_DW01_sub_7n67) );
  XOR2_X2 vscale_core_DW01_sub_7_U67 ( .A(vscale_core_DW01_sub_7n10), .B(vscale_core_DW01_sub_7n73), .Z(pipeline_alu_N272) );
  NAND2_X2 vscale_core_DW01_sub_7_U71 ( .A1(vscale_core_DW01_sub_7n186), .A2(vscale_core_DW01_sub_7n72), .ZN(vscale_core_DW01_sub_7n10) );
  NAND2_X2 vscale_core_DW01_sub_7_U74 ( .A1(vscale_core_DW01_sub_7n217), .A2(pipeline_alu_src_a[19]), .ZN(vscale_core_DW01_sub_7n72) );
  XOR2_X2 vscale_core_DW01_sub_7_U75 ( .A(vscale_core_DW01_sub_7n11), .B(vscale_core_DW01_sub_7n82), .Z(pipeline_alu_N271) );
  NAND2_X2 vscale_core_DW01_sub_7_U79 ( .A1(vscale_core_DW01_sub_7n83), .A2(vscale_core_DW01_sub_7n339), .ZN(vscale_core_DW01_sub_7n76) );
  NAND2_X2 vscale_core_DW01_sub_7_U86 ( .A1(vscale_core_DW01_sub_7n218), .A2(pipeline_alu_src_a[18]), .ZN(vscale_core_DW01_sub_7n81) );
  XOR2_X2 vscale_core_DW01_sub_7_U87 ( .A(vscale_core_DW01_sub_7n12), .B(vscale_core_DW01_sub_7n87), .Z(pipeline_alu_N270) );
  NAND2_X2 vscale_core_DW01_sub_7_U91 ( .A1(vscale_core_DW01_sub_7n188), .A2(vscale_core_DW01_sub_7n86), .ZN(vscale_core_DW01_sub_7n12) );
  XNOR2_X2 vscale_core_DW01_sub_7_U95 ( .A(vscale_core_DW01_sub_7n92), .B(vscale_core_DW01_sub_7n13), .ZN(pipeline_alu_N269) );
  NAND2_X2 vscale_core_DW01_sub_7_U99 ( .A1(vscale_core_DW01_sub_7n88), .A2(vscale_core_DW01_sub_7n91), .ZN(vscale_core_DW01_sub_7n13) );
  XOR2_X2 vscale_core_DW01_sub_7_U103 ( .A(vscale_core_DW01_sub_7n14), .B(vscale_core_DW01_sub_7n102), .Z(pipeline_alu_N268) );
  NAND2_X2 vscale_core_DW01_sub_7_U108 ( .A1(vscale_core_DW01_sub_7n110), .A2(vscale_core_DW01_sub_7n98), .ZN(vscale_core_DW01_sub_7n96) );
  NAND2_X2 vscale_core_DW01_sub_7_U112 ( .A1(vscale_core_DW01_sub_7n190), .A2(vscale_core_DW01_sub_7n101), .ZN(vscale_core_DW01_sub_7n14) );
  XNOR2_X2 vscale_core_DW01_sub_7_U116 ( .A(vscale_core_DW01_sub_7n107), .B(vscale_core_DW01_sub_7n15), .ZN(pipeline_alu_N267) );
  NAND2_X2 vscale_core_DW01_sub_7_U120 ( .A1(vscale_core_DW01_sub_7n191), .A2(vscale_core_DW01_sub_7n106), .ZN(vscale_core_DW01_sub_7n15) );
  NAND2_X2 vscale_core_DW01_sub_7_U123 ( .A1(vscale_core_DW01_sub_7n222), .A2(pipeline_alu_src_a[14]), .ZN(vscale_core_DW01_sub_7n106) );
  XOR2_X2 vscale_core_DW01_sub_7_U124 ( .A(vscale_core_DW01_sub_7n16), .B(vscale_core_DW01_sub_7n114), .Z(pipeline_alu_N266) );
  NAND2_X2 vscale_core_DW01_sub_7_U130 ( .A1(vscale_core_DW01_sub_7n192), .A2(vscale_core_DW01_sub_7n113), .ZN(vscale_core_DW01_sub_7n16) );
  NAND2_X2 vscale_core_DW01_sub_7_U133 ( .A1(vscale_core_DW01_sub_7n223), .A2(n6567), .ZN(vscale_core_DW01_sub_7n113) );
  XOR2_X2 vscale_core_DW01_sub_7_U134 ( .A(vscale_core_DW01_sub_7n17), .B(vscale_core_DW01_sub_7n119), .Z(pipeline_alu_N265) );
  NAND2_X2 vscale_core_DW01_sub_7_U138 ( .A1(vscale_core_DW01_sub_7n193), .A2(vscale_core_DW01_sub_7n118), .ZN(vscale_core_DW01_sub_7n17) );
  XOR2_X2 vscale_core_DW01_sub_7_U142 ( .A(vscale_core_DW01_sub_7n18), .B(vscale_core_DW01_sub_7n127), .Z(pipeline_alu_N264) );
  NAND2_X2 vscale_core_DW01_sub_7_U145 ( .A1(vscale_core_DW01_sub_7n135), .A2(vscale_core_DW01_sub_7n123), .ZN(vscale_core_DW01_sub_7n121) );
  NAND2_X2 vscale_core_DW01_sub_7_U149 ( .A1(vscale_core_DW01_sub_7n194), .A2(vscale_core_DW01_sub_7n126), .ZN(vscale_core_DW01_sub_7n18) );
  XNOR2_X2 vscale_core_DW01_sub_7_U153 ( .A(vscale_core_DW01_sub_7n132), .B(vscale_core_DW01_sub_7n19), .ZN(pipeline_alu_N263) );
  NAND2_X2 vscale_core_DW01_sub_7_U157 ( .A1(vscale_core_DW01_sub_7n195), .A2(vscale_core_DW01_sub_7n131), .ZN(vscale_core_DW01_sub_7n19) );
  XNOR2_X2 vscale_core_DW01_sub_7_U161 ( .A(vscale_core_DW01_sub_7n139), .B(vscale_core_DW01_sub_7n20), .ZN(pipeline_alu_N262) );
  NAND2_X2 vscale_core_DW01_sub_7_U167 ( .A1(vscale_core_DW01_sub_7n196), .A2(vscale_core_DW01_sub_7n138), .ZN(vscale_core_DW01_sub_7n20) );
  NAND2_X2 vscale_core_DW01_sub_7_U170 ( .A1(vscale_core_DW01_sub_7n227), .A2(n6973), .ZN(vscale_core_DW01_sub_7n138) );
  XOR2_X2 vscale_core_DW01_sub_7_U171 ( .A(vscale_core_DW01_sub_7n21), .B(vscale_core_DW01_sub_7n142), .Z(pipeline_alu_N261) );
  NAND2_X2 vscale_core_DW01_sub_7_U173 ( .A1(vscale_core_DW01_sub_7n197), .A2(vscale_core_DW01_sub_7n141), .ZN(vscale_core_DW01_sub_7n21) );
  XNOR2_X2 vscale_core_DW01_sub_7_U177 ( .A(vscale_core_DW01_sub_7n150), .B(vscale_core_DW01_sub_7n22), .ZN(pipeline_alu_N260) );
  NAND2_X2 vscale_core_DW01_sub_7_U180 ( .A1(vscale_core_DW01_sub_7n154), .A2(vscale_core_DW01_sub_7n146), .ZN(vscale_core_DW01_sub_7n144) );
  XOR2_X2 vscale_core_DW01_sub_7_U188 ( .A(vscale_core_DW01_sub_7n23), .B(vscale_core_DW01_sub_7n153), .Z(pipeline_alu_N259) );
  NAND2_X2 vscale_core_DW01_sub_7_U190 ( .A1(vscale_core_DW01_sub_7n199), .A2(vscale_core_DW01_sub_7n152), .ZN(vscale_core_DW01_sub_7n23) );
  XOR2_X2 vscale_core_DW01_sub_7_U194 ( .A(vscale_core_DW01_sub_7n24), .B(vscale_core_DW01_sub_7n158), .Z(pipeline_alu_N258) );
  XNOR2_X2 vscale_core_DW01_sub_7_U202 ( .A(vscale_core_DW01_sub_7n163), .B(vscale_core_DW01_sub_7n25), .ZN(pipeline_alu_N257) );
  XNOR2_X2 vscale_core_DW01_sub_7_U210 ( .A(vscale_core_DW01_sub_7n169), .B(vscale_core_DW01_sub_7n26), .ZN(pipeline_alu_N256) );
  NAND2_X2 vscale_core_DW01_sub_7_U215 ( .A1(vscale_core_DW01_sub_7n202), .A2(vscale_core_DW01_sub_7n168), .ZN(vscale_core_DW01_sub_7n26) );
  NAND2_X2 vscale_core_DW01_sub_7_U218 ( .A1(vscale_core_DW01_sub_7n233), .A2(n6634), .ZN(vscale_core_DW01_sub_7n168) );
  XOR2_X2 vscale_core_DW01_sub_7_U219 ( .A(vscale_core_DW01_sub_7n27), .B(vscale_core_DW01_sub_7n172), .Z(pipeline_alu_N255) );
  NAND2_X2 vscale_core_DW01_sub_7_U221 ( .A1(vscale_core_DW01_sub_7n203), .A2(vscale_core_DW01_sub_7n171), .ZN(vscale_core_DW01_sub_7n27) );
  NAND2_X2 vscale_core_DW01_sub_7_U231 ( .A1(vscale_core_DW01_sub_7n235), .A2(n6632), .ZN(vscale_core_DW01_sub_7n175) );
  INV_X1 vscale_core_DW01_sub_7_U269 ( .A(pipeline_alu_src_b[8]), .ZN(vscale_core_DW01_sub_7n228) );
  AOI21_X2 vscale_core_DW01_sub_7_U270 ( .B1(vscale_core_DW01_sub_7n61), .B2(vscale_core_DW01_sub_7n341), .A(vscale_core_DW01_sub_7n58), .ZN(vscale_core_DW01_sub_7n56) );
  OAI21_X2 vscale_core_DW01_sub_7_U271 ( .B1(vscale_core_DW01_sub_7n56), .B2(vscale_core_DW01_sub_7n54), .A(vscale_core_DW01_sub_7n55), .ZN(vscale_core_DW01_sub_7n53) );
  AOI21_X2 vscale_core_DW01_sub_7_U272 ( .B1(vscale_core_DW01_sub_7n45), .B2(vscale_core_DW01_sub_7n344), .A(vscale_core_DW01_sub_7n42), .ZN(vscale_core_DW01_sub_7n40) );
  INV_X1 vscale_core_DW01_sub_7_U273 ( .A(pipeline_alu_src_b[7]), .ZN(vscale_core_DW01_sub_7n229) );
  OAI21_X2 vscale_core_DW01_sub_7_U274 ( .B1(vscale_core_DW01_sub_7n93), .B2(vscale_core_DW01_sub_7n62), .A(vscale_core_DW01_sub_7n63), .ZN(vscale_core_DW01_sub_7n61) );
  AOI21_X2 vscale_core_DW01_sub_7_U275 ( .B1(vscale_core_DW01_sub_7n53), .B2(vscale_core_DW01_sub_7n342), .A(vscale_core_DW01_sub_7n50), .ZN(vscale_core_DW01_sub_7n48) );
  OAI21_X2 vscale_core_DW01_sub_7_U276 ( .B1(vscale_core_DW01_sub_7n48), .B2(vscale_core_DW01_sub_7n46), .A(vscale_core_DW01_sub_7n47), .ZN(vscale_core_DW01_sub_7n45) );
  INV_X1 vscale_core_DW01_sub_7_U277 ( .A(n6556), .ZN(vscale_core_DW01_sub_7n207) );
  INV_X1 vscale_core_DW01_sub_7_U278 ( .A(pipeline_alu_src_b[28]), .ZN(vscale_core_DW01_sub_7n208) );
  INV_X1 vscale_core_DW01_sub_7_U279 ( .A(pipeline_alu_src_b[12]), .ZN(vscale_core_DW01_sub_7n224) );
  INV_X2 vscale_core_DW01_sub_7_U280 ( .A(pipeline_alu_src_b[16]), .ZN(vscale_core_DW01_sub_7n220) );
  INV_X1 vscale_core_DW01_sub_7_U281 ( .A(pipeline_alu_src_b[15]), .ZN(vscale_core_DW01_sub_7n221) );
  AOI21_X4 vscale_core_DW01_sub_7_U282 ( .B1(vscale_core_DW01_sub_7n143), .B2(vscale_core_DW01_sub_7n94), .A(vscale_core_DW01_sub_7n95), .ZN(vscale_core_DW01_sub_7n93) );
  INV_X2 vscale_core_DW01_sub_7_U283 ( .A(pipeline_alu_src_b[21]), .ZN(vscale_core_DW01_sub_7n215) );
  NAND2_X1 vscale_core_DW01_sub_7_U284 ( .A1(vscale_core_DW01_sub_7n229), .A2(n6611), .ZN(vscale_core_DW01_sub_7n149) );
  NAND2_X1 vscale_core_DW01_sub_7_U285 ( .A1(vscale_core_DW01_sub_7n231), .A2(n6621), .ZN(vscale_core_DW01_sub_7n157) );
  NAND2_X1 vscale_core_DW01_sub_7_U286 ( .A1(vscale_core_DW01_sub_7n234), .A2(pipeline_alu_src_a[2]), .ZN(vscale_core_DW01_sub_7n171) );
  XNOR2_X1 vscale_core_DW01_sub_7_U287 ( .A(vscale_core_DW01_sub_7n236), .B(pipeline_alu_src_a[0]), .ZN(pipeline_alu_N253) );
  INV_X2 vscale_core_DW01_sub_7_U288 ( .A(pipeline_alu_src_b[5]), .ZN(vscale_core_DW01_sub_7n231) );
  NAND2_X1 vscale_core_DW01_sub_7_U289 ( .A1(vscale_core_DW01_sub_7n225), .A2(n6614), .ZN(vscale_core_DW01_sub_7n126) );
  NAND2_X1 vscale_core_DW01_sub_7_U290 ( .A1(vscale_core_DW01_sub_7n209), .A2(n6602), .ZN(vscale_core_DW01_sub_7n36) );
  NAND2_X1 vscale_core_DW01_sub_7_U291 ( .A1(vscale_core_DW01_sub_7n219), .A2(pipeline_alu_src_a[17]), .ZN(vscale_core_DW01_sub_7n86) );
  NAND2_X1 vscale_core_DW01_sub_7_U292 ( .A1(vscale_core_DW01_sub_7n232), .A2(n6927), .ZN(vscale_core_DW01_sub_7n162) );
  NOR2_X1 vscale_core_DW01_sub_7_U293 ( .A1(vscale_core_DW01_sub_7n170), .A2(vscale_core_DW01_sub_7n167), .ZN(vscale_core_DW01_sub_7n165) );
  OAI21_X1 vscale_core_DW01_sub_7_U294 ( .B1(vscale_core_DW01_sub_7n112), .B2(vscale_core_DW01_sub_7n118), .A(vscale_core_DW01_sub_7n113), .ZN(vscale_core_DW01_sub_7n111) );
  OAI21_X1 vscale_core_DW01_sub_7_U295 ( .B1(vscale_core_DW01_sub_7n85), .B2(vscale_core_DW01_sub_7n91), .A(vscale_core_DW01_sub_7n86), .ZN(vscale_core_DW01_sub_7n84) );
  NOR2_X1 vscale_core_DW01_sub_7_U296 ( .A1(vscale_core_DW01_sub_7n117), .A2(vscale_core_DW01_sub_7n112), .ZN(vscale_core_DW01_sub_7n110) );
  NAND2_X1 vscale_core_DW01_sub_7_U297 ( .A1(vscale_core_DW01_sub_7n201), .A2(vscale_core_DW01_sub_7n162), .ZN(vscale_core_DW01_sub_7n25) );
  INV_X1 vscale_core_DW01_sub_7_U298 ( .A(vscale_core_DW01_sub_7n161), .ZN(vscale_core_DW01_sub_7n201) );
  OAI21_X1 vscale_core_DW01_sub_7_U299 ( .B1(vscale_core_DW01_sub_7n142), .B2(vscale_core_DW01_sub_7n140), .A(vscale_core_DW01_sub_7n141), .ZN(vscale_core_DW01_sub_7n139) );
  NOR2_X2 vscale_core_DW01_sub_7_U300 ( .A1(vscale_core_DW01_sub_7n76), .A2(vscale_core_DW01_sub_7n71), .ZN(vscale_core_DW01_sub_7n69) );
  AOI21_X1 vscale_core_DW01_sub_7_U301 ( .B1(vscale_core_DW01_sub_7n163), .B2(vscale_core_DW01_sub_7n154), .A(vscale_core_DW01_sub_7n155), .ZN(vscale_core_DW01_sub_7n153) );
  OAI21_X1 vscale_core_DW01_sub_7_U302 ( .B1(vscale_core_DW01_sub_7n142), .B2(vscale_core_DW01_sub_7n121), .A(vscale_core_DW01_sub_7n122), .ZN(vscale_core_DW01_sub_7n120) );
  INV_X1 vscale_core_DW01_sub_7_U303 ( .A(vscale_core_DW01_sub_7n173), .ZN(vscale_core_DW01_sub_7n172) );
  OAI21_X1 vscale_core_DW01_sub_7_U304 ( .B1(vscale_core_DW01_sub_7n167), .B2(vscale_core_DW01_sub_7n171), .A(vscale_core_DW01_sub_7n168), .ZN(vscale_core_DW01_sub_7n166) );
  OAI21_X1 vscale_core_DW01_sub_7_U305 ( .B1(vscale_core_DW01_sub_7n137), .B2(vscale_core_DW01_sub_7n141), .A(vscale_core_DW01_sub_7n138), .ZN(vscale_core_DW01_sub_7n136) );
  NOR2_X1 vscale_core_DW01_sub_7_U306 ( .A1(vscale_core_DW01_sub_7n140), .A2(vscale_core_DW01_sub_7n137), .ZN(vscale_core_DW01_sub_7n135) );
  OAI21_X1 vscale_core_DW01_sub_7_U307 ( .B1(vscale_core_DW01_sub_7n148), .B2(vscale_core_DW01_sub_7n152), .A(vscale_core_DW01_sub_7n149), .ZN(vscale_core_DW01_sub_7n147) );
  NOR2_X1 vscale_core_DW01_sub_7_U308 ( .A1(vscale_core_DW01_sub_7n161), .A2(vscale_core_DW01_sub_7n156), .ZN(vscale_core_DW01_sub_7n154) );
  NOR2_X1 vscale_core_DW01_sub_7_U309 ( .A1(vscale_core_DW01_sub_7n130), .A2(vscale_core_DW01_sub_7n125), .ZN(vscale_core_DW01_sub_7n123) );
  NOR2_X1 vscale_core_DW01_sub_7_U310 ( .A1(vscale_core_DW01_sub_7n85), .A2(vscale_core_DW01_sub_7n90), .ZN(vscale_core_DW01_sub_7n83) );
  NAND2_X1 vscale_core_DW01_sub_7_U311 ( .A1(vscale_core_DW01_sub_7n339), .A2(vscale_core_DW01_sub_7n81), .ZN(vscale_core_DW01_sub_7n11) );
  INV_X1 vscale_core_DW01_sub_7_U312 ( .A(vscale_core_DW01_sub_7n100), .ZN(vscale_core_DW01_sub_7n190) );
  INV_X1 vscale_core_DW01_sub_7_U313 ( .A(vscale_core_DW01_sub_7n85), .ZN(vscale_core_DW01_sub_7n188) );
  INV_X1 vscale_core_DW01_sub_7_U314 ( .A(vscale_core_DW01_sub_7n71), .ZN(vscale_core_DW01_sub_7n186) );
  XOR2_X1 vscale_core_DW01_sub_7_U315 ( .A(vscale_core_DW01_sub_7n176), .B(vscale_core_DW01_sub_7n28), .Z(pipeline_alu_N254) );
  NAND2_X1 vscale_core_DW01_sub_7_U316 ( .A1(vscale_core_DW01_sub_7n204), .A2(vscale_core_DW01_sub_7n175), .ZN(vscale_core_DW01_sub_7n28) );
  INV_X1 vscale_core_DW01_sub_7_U317 ( .A(vscale_core_DW01_sub_7n174), .ZN(vscale_core_DW01_sub_7n204) );
  OAI21_X1 vscale_core_DW01_sub_7_U318 ( .B1(vscale_core_DW01_sub_7n172), .B2(vscale_core_DW01_sub_7n170), .A(vscale_core_DW01_sub_7n171), .ZN(vscale_core_DW01_sub_7n169) );
  INV_X1 vscale_core_DW01_sub_7_U319 ( .A(vscale_core_DW01_sub_7n167), .ZN(vscale_core_DW01_sub_7n202) );
  NAND2_X1 vscale_core_DW01_sub_7_U320 ( .A1(vscale_core_DW01_sub_7n200), .A2(vscale_core_DW01_sub_7n157), .ZN(vscale_core_DW01_sub_7n24) );
  INV_X1 vscale_core_DW01_sub_7_U321 ( .A(vscale_core_DW01_sub_7n156), .ZN(vscale_core_DW01_sub_7n200) );
  NAND2_X1 vscale_core_DW01_sub_7_U322 ( .A1(vscale_core_DW01_sub_7n198), .A2(vscale_core_DW01_sub_7n149), .ZN(vscale_core_DW01_sub_7n22) );
  INV_X1 vscale_core_DW01_sub_7_U323 ( .A(vscale_core_DW01_sub_7n148), .ZN(vscale_core_DW01_sub_7n198) );
  XNOR2_X1 vscale_core_DW01_sub_7_U324 ( .A(n7005), .B(n13159), .ZN(vscale_core_DW01_sub_7n1) );
  NOR2_X2 vscale_core_DW01_sub_7_U325 ( .A1(vscale_core_DW01_sub_7n121), .A2(vscale_core_DW01_sub_7n96), .ZN(vscale_core_DW01_sub_7n94) );
  OAI21_X2 vscale_core_DW01_sub_7_U326 ( .B1(vscale_core_DW01_sub_7n122), .B2(vscale_core_DW01_sub_7n96), .A(vscale_core_DW01_sub_7n97), .ZN(vscale_core_DW01_sub_7n95) );
  OAI21_X2 vscale_core_DW01_sub_7_U327 ( .B1(vscale_core_DW01_sub_7n142), .B2(vscale_core_DW01_sub_7n133), .A(vscale_core_DW01_sub_7n134), .ZN(vscale_core_DW01_sub_7n132) );
  OAI21_X2 vscale_core_DW01_sub_7_U328 ( .B1(vscale_core_DW01_sub_7n119), .B2(vscale_core_DW01_sub_7n108), .A(vscale_core_DW01_sub_7n109), .ZN(vscale_core_DW01_sub_7n107) );
  AOI21_X2 vscale_core_DW01_sub_7_U329 ( .B1(vscale_core_DW01_sub_7n123), .B2(vscale_core_DW01_sub_7n136), .A(vscale_core_DW01_sub_7n124), .ZN(vscale_core_DW01_sub_7n122) );
  OAI21_X1 vscale_core_DW01_sub_7_U330 ( .B1(vscale_core_DW01_sub_7n125), .B2(vscale_core_DW01_sub_7n131), .A(vscale_core_DW01_sub_7n126), .ZN(vscale_core_DW01_sub_7n124) );
  AOI21_X2 vscale_core_DW01_sub_7_U331 ( .B1(vscale_core_DW01_sub_7n84), .B2(vscale_core_DW01_sub_7n339), .A(vscale_core_DW01_sub_7n79), .ZN(vscale_core_DW01_sub_7n77) );
  AOI21_X2 vscale_core_DW01_sub_7_U332 ( .B1(vscale_core_DW01_sub_7n165), .B2(vscale_core_DW01_sub_7n173), .A(vscale_core_DW01_sub_7n166), .ZN(vscale_core_DW01_sub_7n164) );
  OAI21_X2 vscale_core_DW01_sub_7_U333 ( .B1(vscale_core_DW01_sub_7n156), .B2(vscale_core_DW01_sub_7n162), .A(vscale_core_DW01_sub_7n157), .ZN(vscale_core_DW01_sub_7n155) );
  OAI21_X2 vscale_core_DW01_sub_7_U334 ( .B1(vscale_core_DW01_sub_7n77), .B2(vscale_core_DW01_sub_7n71), .A(vscale_core_DW01_sub_7n72), .ZN(vscale_core_DW01_sub_7n70) );
  OAI21_X2 vscale_core_DW01_sub_7_U335 ( .B1(vscale_core_DW01_sub_7n40), .B2(vscale_core_DW01_sub_7n38), .A(vscale_core_DW01_sub_7n39), .ZN(vscale_core_DW01_sub_7n37) );
  AOI21_X2 vscale_core_DW01_sub_7_U336 ( .B1(vscale_core_DW01_sub_7n70), .B2(vscale_core_DW01_sub_7n340), .A(vscale_core_DW01_sub_7n65), .ZN(vscale_core_DW01_sub_7n63) );
  OAI21_X2 vscale_core_DW01_sub_7_U337 ( .B1(vscale_core_DW01_sub_7n174), .B2(vscale_core_DW01_sub_7n176), .A(vscale_core_DW01_sub_7n175), .ZN(vscale_core_DW01_sub_7n173) );
  AOI21_X2 vscale_core_DW01_sub_7_U338 ( .B1(vscale_core_DW01_sub_7n98), .B2(vscale_core_DW01_sub_7n111), .A(vscale_core_DW01_sub_7n99), .ZN(vscale_core_DW01_sub_7n97) );
  OAI21_X1 vscale_core_DW01_sub_7_U339 ( .B1(vscale_core_DW01_sub_7n100), .B2(vscale_core_DW01_sub_7n106), .A(vscale_core_DW01_sub_7n101), .ZN(vscale_core_DW01_sub_7n99) );
  OAI21_X2 vscale_core_DW01_sub_7_U340 ( .B1(vscale_core_DW01_sub_7n164), .B2(vscale_core_DW01_sub_7n144), .A(vscale_core_DW01_sub_7n145), .ZN(vscale_core_DW01_sub_7n143) );
  AOI21_X2 vscale_core_DW01_sub_7_U341 ( .B1(vscale_core_DW01_sub_7n155), .B2(vscale_core_DW01_sub_7n146), .A(vscale_core_DW01_sub_7n147), .ZN(vscale_core_DW01_sub_7n145) );
  NOR2_X2 vscale_core_DW01_sub_7_U342 ( .A1(vscale_core_DW01_sub_7n151), .A2(vscale_core_DW01_sub_7n148), .ZN(vscale_core_DW01_sub_7n146) );
  NOR2_X1 vscale_core_DW01_sub_7_U343 ( .A1(vscale_core_DW01_sub_7n105), .A2(vscale_core_DW01_sub_7n100), .ZN(vscale_core_DW01_sub_7n98) );
  AOI21_X2 vscale_core_DW01_sub_7_U344 ( .B1(vscale_core_DW01_sub_7n107), .B2(vscale_core_DW01_sub_7n191), .A(vscale_core_DW01_sub_7n104), .ZN(vscale_core_DW01_sub_7n102) );
  AOI21_X2 vscale_core_DW01_sub_7_U345 ( .B1(vscale_core_DW01_sub_7n92), .B2(vscale_core_DW01_sub_7n88), .A(vscale_core_DW01_sub_7n89), .ZN(vscale_core_DW01_sub_7n87) );
  AOI21_X1 vscale_core_DW01_sub_7_U346 ( .B1(vscale_core_DW01_sub_7n92), .B2(vscale_core_DW01_sub_7n83), .A(vscale_core_DW01_sub_7n84), .ZN(vscale_core_DW01_sub_7n82) );
  AOI21_X2 vscale_core_DW01_sub_7_U347 ( .B1(vscale_core_DW01_sub_7n92), .B2(vscale_core_DW01_sub_7n74), .A(vscale_core_DW01_sub_7n75), .ZN(vscale_core_DW01_sub_7n73) );
  AOI21_X1 vscale_core_DW01_sub_7_U348 ( .B1(vscale_core_DW01_sub_7n92), .B2(vscale_core_DW01_sub_7n69), .A(vscale_core_DW01_sub_7n70), .ZN(vscale_core_DW01_sub_7n68) );
  AOI21_X2 vscale_core_DW01_sub_7_U349 ( .B1(vscale_core_DW01_sub_7n132), .B2(vscale_core_DW01_sub_7n195), .A(vscale_core_DW01_sub_7n129), .ZN(vscale_core_DW01_sub_7n127) );
  AOI21_X2 vscale_core_DW01_sub_7_U350 ( .B1(vscale_core_DW01_sub_7n120), .B2(vscale_core_DW01_sub_7n193), .A(vscale_core_DW01_sub_7n116), .ZN(vscale_core_DW01_sub_7n114) );
  OAI21_X1 vscale_core_DW01_sub_7_U351 ( .B1(vscale_core_DW01_sub_7n153), .B2(vscale_core_DW01_sub_7n151), .A(vscale_core_DW01_sub_7n152), .ZN(vscale_core_DW01_sub_7n150) );
  AOI21_X2 vscale_core_DW01_sub_7_U352 ( .B1(vscale_core_DW01_sub_7n163), .B2(vscale_core_DW01_sub_7n201), .A(vscale_core_DW01_sub_7n160), .ZN(vscale_core_DW01_sub_7n158) );
  NOR2_X1 vscale_core_DW01_sub_7_U353 ( .A1(vscale_core_DW01_sub_7n219), .A2(pipeline_alu_src_a[17]), .ZN(vscale_core_DW01_sub_7n85) );
  NOR2_X1 vscale_core_DW01_sub_7_U354 ( .A1(vscale_core_DW01_sub_7n233), .A2(n6634), .ZN(vscale_core_DW01_sub_7n167) );
  NOR2_X1 vscale_core_DW01_sub_7_U355 ( .A1(vscale_core_DW01_sub_7n223), .A2(n6567), .ZN(vscale_core_DW01_sub_7n112) );
  NOR2_X1 vscale_core_DW01_sub_7_U356 ( .A1(vscale_core_DW01_sub_7n225), .A2(n6614), .ZN(vscale_core_DW01_sub_7n125) );
  NOR2_X1 vscale_core_DW01_sub_7_U357 ( .A1(vscale_core_DW01_sub_7n227), .A2(n6973), .ZN(vscale_core_DW01_sub_7n137) );
  NOR2_X1 vscale_core_DW01_sub_7_U358 ( .A1(vscale_core_DW01_sub_7n229), .A2(n6611), .ZN(vscale_core_DW01_sub_7n148) );
  NOR2_X1 vscale_core_DW01_sub_7_U359 ( .A1(vscale_core_DW01_sub_7n231), .A2(n6621), .ZN(vscale_core_DW01_sub_7n156) );
  AOI21_X2 vscale_core_DW01_sub_7_U360 ( .B1(vscale_core_DW01_sub_7n37), .B2(vscale_core_DW01_sub_7n343), .A(vscale_core_DW01_sub_7n34), .ZN(vscale_core_DW01_sub_7n32) );
  NOR2_X1 vscale_core_DW01_sub_7_U361 ( .A1(vscale_core_DW01_sub_7n234), .A2(pipeline_alu_src_a[2]), .ZN(vscale_core_DW01_sub_7n170) );
  NOR2_X1 vscale_core_DW01_sub_7_U362 ( .A1(vscale_core_DW01_sub_7n217), .A2(pipeline_alu_src_a[19]), .ZN(vscale_core_DW01_sub_7n71) );
  NOR2_X1 vscale_core_DW01_sub_7_U363 ( .A1(vscale_core_DW01_sub_7n214), .A2(n6625), .ZN(vscale_core_DW01_sub_7n54) );
  NOR2_X1 vscale_core_DW01_sub_7_U364 ( .A1(vscale_core_DW01_sub_7n235), .A2(n6632), .ZN(vscale_core_DW01_sub_7n174) );
  NOR2_X1 vscale_core_DW01_sub_7_U365 ( .A1(vscale_core_DW01_sub_7n232), .A2(n6927), .ZN(vscale_core_DW01_sub_7n161) );
  NOR2_X1 vscale_core_DW01_sub_7_U366 ( .A1(vscale_core_DW01_sub_7n222), .A2(pipeline_alu_src_a[14]), .ZN(vscale_core_DW01_sub_7n105) );
  NOR2_X1 vscale_core_DW01_sub_7_U367 ( .A1(vscale_core_DW01_sub_7n236), .A2(pipeline_alu_src_a[0]), .ZN(vscale_core_DW01_sub_7n176) );
  OR2_X1 vscale_core_DW01_sub_7_U368 ( .A1(vscale_core_DW01_sub_7n218), .A2(pipeline_alu_src_a[18]), .ZN(vscale_core_DW01_sub_7n339) );
  OR2_X1 vscale_core_DW01_sub_7_U369 ( .A1(vscale_core_DW01_sub_7n216), .A2(pipeline_alu_src_a[20]), .ZN(vscale_core_DW01_sub_7n340) );
  OR2_X1 vscale_core_DW01_sub_7_U370 ( .A1(vscale_core_DW01_sub_7n215), .A2(pipeline_alu_src_a[21]), .ZN(vscale_core_DW01_sub_7n341) );
  NOR2_X1 vscale_core_DW01_sub_7_U371 ( .A1(vscale_core_DW01_sub_7n212), .A2(pipeline_alu_src_a[24]), .ZN(vscale_core_DW01_sub_7n46) );
  NOR2_X1 vscale_core_DW01_sub_7_U372 ( .A1(vscale_core_DW01_sub_7n210), .A2(n6561), .ZN(vscale_core_DW01_sub_7n38) );
  OR2_X1 vscale_core_DW01_sub_7_U373 ( .A1(vscale_core_DW01_sub_7n213), .A2(n6980), .ZN(vscale_core_DW01_sub_7n342) );
  OR2_X1 vscale_core_DW01_sub_7_U374 ( .A1(vscale_core_DW01_sub_7n209), .A2(n6602), .ZN(vscale_core_DW01_sub_7n343) );
  OR2_X1 vscale_core_DW01_sub_7_U375 ( .A1(vscale_core_DW01_sub_7n211), .A2(n6609), .ZN(vscale_core_DW01_sub_7n344) );
  INV_X1 vscale_core_DW01_sub_7_U376 ( .A(pipeline_alu_src_b[27]), .ZN(vscale_core_DW01_sub_7n209) );
  NOR2_X1 vscale_core_DW01_sub_7_U377 ( .A1(vscale_core_DW01_sub_7n226), .A2(n6572), .ZN(vscale_core_DW01_sub_7n130) );
  NAND2_X1 vscale_core_DW01_sub_7_U378 ( .A1(vscale_core_DW01_sub_7n226), .A2(n6572), .ZN(vscale_core_DW01_sub_7n131) );
  INV_X2 vscale_core_DW01_sub_7_U379 ( .A(pipeline_alu_src_b[14]), .ZN(vscale_core_DW01_sub_7n222) );
  NOR2_X1 vscale_core_DW01_sub_7_U380 ( .A1(vscale_core_DW01_sub_7n224), .A2(pipeline_alu_src_a[12]), .ZN(vscale_core_DW01_sub_7n117) );
  NAND2_X1 vscale_core_DW01_sub_7_U381 ( .A1(vscale_core_DW01_sub_7n224), .A2(pipeline_alu_src_a[12]), .ZN(vscale_core_DW01_sub_7n118) );
  INV_X2 vscale_core_DW01_sub_7_U382 ( .A(n6976), .ZN(vscale_core_DW01_sub_7n235) );
  NAND2_X1 vscale_core_DW01_sub_7_U383 ( .A1(vscale_core_DW01_sub_7n221), .A2(n6597), .ZN(vscale_core_DW01_sub_7n101) );
  NOR2_X1 vscale_core_DW01_sub_7_U384 ( .A1(vscale_core_DW01_sub_7n221), .A2(n6597), .ZN(vscale_core_DW01_sub_7n100) );
  NOR2_X1 vscale_core_DW01_sub_7_U385 ( .A1(vscale_core_DW01_sub_7n220), .A2(pipeline_alu_src_a[16]), .ZN(vscale_core_DW01_sub_7n90) );
  NAND2_X1 vscale_core_DW01_sub_7_U386 ( .A1(vscale_core_DW01_sub_7n220), .A2(pipeline_alu_src_a[16]), .ZN(vscale_core_DW01_sub_7n91) );
  NOR2_X1 vscale_core_DW01_sub_7_U387 ( .A1(vscale_core_DW01_sub_7n230), .A2(n6605), .ZN(vscale_core_DW01_sub_7n151) );
  NAND2_X1 vscale_core_DW01_sub_7_U388 ( .A1(vscale_core_DW01_sub_7n230), .A2(n6605), .ZN(vscale_core_DW01_sub_7n152) );
  NOR2_X1 vscale_core_DW01_sub_7_U389 ( .A1(vscale_core_DW01_sub_7n228), .A2(n9335), .ZN(vscale_core_DW01_sub_7n140) );
  NAND2_X1 vscale_core_DW01_sub_7_U390 ( .A1(vscale_core_DW01_sub_7n228), .A2(n9335), .ZN(vscale_core_DW01_sub_7n141) );
  INV_X2 vscale_core_DW01_sub_7_U391 ( .A(n9339), .ZN(vscale_core_DW01_sub_7n233) );
  INV_X4 vscale_core_DW01_sub_7_U392 ( .A(vscale_core_DW01_sub_7n93), .ZN(vscale_core_DW01_sub_7n92) );
  INV_X4 vscale_core_DW01_sub_7_U393 ( .A(vscale_core_DW01_sub_7n91), .ZN(vscale_core_DW01_sub_7n89) );
  INV_X4 vscale_core_DW01_sub_7_U394 ( .A(vscale_core_DW01_sub_7n81), .ZN(vscale_core_DW01_sub_7n79) );
  INV_X4 vscale_core_DW01_sub_7_U395 ( .A(vscale_core_DW01_sub_7n77), .ZN(vscale_core_DW01_sub_7n75) );
  INV_X4 vscale_core_DW01_sub_7_U396 ( .A(vscale_core_DW01_sub_7n76), .ZN(vscale_core_DW01_sub_7n74) );
  INV_X4 vscale_core_DW01_sub_7_U397 ( .A(vscale_core_DW01_sub_7n67), .ZN(vscale_core_DW01_sub_7n65) );
  INV_X4 vscale_core_DW01_sub_7_U398 ( .A(vscale_core_DW01_sub_7n60), .ZN(vscale_core_DW01_sub_7n58) );
  INV_X4 vscale_core_DW01_sub_7_U399 ( .A(vscale_core_DW01_sub_7n52), .ZN(vscale_core_DW01_sub_7n50) );
  INV_X4 vscale_core_DW01_sub_7_U400 ( .A(vscale_core_DW01_sub_7n44), .ZN(vscale_core_DW01_sub_7n42) );
  INV_X4 vscale_core_DW01_sub_7_U401 ( .A(vscale_core_DW01_sub_7n36), .ZN(vscale_core_DW01_sub_7n34) );
  INV_X4 vscale_core_DW01_sub_7_U402 ( .A(n6617), .ZN(vscale_core_DW01_sub_7n236) );
  INV_X4 vscale_core_DW01_sub_7_U403 ( .A(n9398), .ZN(vscale_core_DW01_sub_7n234) );
  INV_X4 vscale_core_DW01_sub_7_U404 ( .A(pipeline_alu_src_b[4]), .ZN(vscale_core_DW01_sub_7n232) );
  INV_X4 vscale_core_DW01_sub_7_U405 ( .A(pipeline_alu_src_b[6]), .ZN(vscale_core_DW01_sub_7n230) );
  INV_X4 vscale_core_DW01_sub_7_U406 ( .A(pipeline_alu_src_b[9]), .ZN(vscale_core_DW01_sub_7n227) );
  INV_X4 vscale_core_DW01_sub_7_U407 ( .A(pipeline_alu_src_b[10]), .ZN(vscale_core_DW01_sub_7n226) );
  INV_X4 vscale_core_DW01_sub_7_U408 ( .A(pipeline_alu_src_b[11]), .ZN(vscale_core_DW01_sub_7n225) );
  INV_X4 vscale_core_DW01_sub_7_U409 ( .A(pipeline_alu_src_b[13]), .ZN(vscale_core_DW01_sub_7n223) );
  INV_X4 vscale_core_DW01_sub_7_U410 ( .A(pipeline_alu_src_b[17]), .ZN(vscale_core_DW01_sub_7n219) );
  INV_X4 vscale_core_DW01_sub_7_U411 ( .A(pipeline_alu_src_b[18]), .ZN(vscale_core_DW01_sub_7n218) );
  INV_X4 vscale_core_DW01_sub_7_U412 ( .A(pipeline_alu_src_b[19]), .ZN(vscale_core_DW01_sub_7n217) );
  INV_X4 vscale_core_DW01_sub_7_U413 ( .A(pipeline_alu_src_b[20]), .ZN(vscale_core_DW01_sub_7n216) );
  INV_X4 vscale_core_DW01_sub_7_U414 ( .A(pipeline_alu_src_b[22]), .ZN(vscale_core_DW01_sub_7n214) );
  INV_X4 vscale_core_DW01_sub_7_U415 ( .A(pipeline_alu_src_b[23]), .ZN(vscale_core_DW01_sub_7n213) );
  INV_X4 vscale_core_DW01_sub_7_U416 ( .A(pipeline_alu_src_b[24]), .ZN(vscale_core_DW01_sub_7n212) );
  INV_X4 vscale_core_DW01_sub_7_U417 ( .A(pipeline_alu_src_b[25]), .ZN(vscale_core_DW01_sub_7n211) );
  INV_X4 vscale_core_DW01_sub_7_U418 ( .A(pipeline_alu_src_b[26]), .ZN(vscale_core_DW01_sub_7n210) );
  INV_X4 vscale_core_DW01_sub_7_U419 ( .A(pipeline_alu_src_b[30]), .ZN(vscale_core_DW01_sub_7n206) );
  INV_X4 vscale_core_DW01_sub_7_U420 ( .A(vscale_core_DW01_sub_7n170), .ZN(vscale_core_DW01_sub_7n203) );
  INV_X4 vscale_core_DW01_sub_7_U421 ( .A(vscale_core_DW01_sub_7n151), .ZN(vscale_core_DW01_sub_7n199) );
  INV_X4 vscale_core_DW01_sub_7_U422 ( .A(vscale_core_DW01_sub_7n140), .ZN(vscale_core_DW01_sub_7n197) );
  INV_X4 vscale_core_DW01_sub_7_U423 ( .A(vscale_core_DW01_sub_7n137), .ZN(vscale_core_DW01_sub_7n196) );
  INV_X4 vscale_core_DW01_sub_7_U424 ( .A(vscale_core_DW01_sub_7n125), .ZN(vscale_core_DW01_sub_7n194) );
  INV_X4 vscale_core_DW01_sub_7_U425 ( .A(vscale_core_DW01_sub_7n112), .ZN(vscale_core_DW01_sub_7n192) );
  INV_X4 vscale_core_DW01_sub_7_U426 ( .A(vscale_core_DW01_sub_7n90), .ZN(vscale_core_DW01_sub_7n88) );
  INV_X4 vscale_core_DW01_sub_7_U427 ( .A(vscale_core_DW01_sub_7n54), .ZN(vscale_core_DW01_sub_7n183) );
  INV_X4 vscale_core_DW01_sub_7_U428 ( .A(vscale_core_DW01_sub_7n46), .ZN(vscale_core_DW01_sub_7n181) );
  INV_X4 vscale_core_DW01_sub_7_U429 ( .A(vscale_core_DW01_sub_7n38), .ZN(vscale_core_DW01_sub_7n179) );
  INV_X4 vscale_core_DW01_sub_7_U430 ( .A(vscale_core_DW01_sub_7n32), .ZN(vscale_core_DW01_sub_7n177) );
  INV_X4 vscale_core_DW01_sub_7_U431 ( .A(vscale_core_DW01_sub_7n164), .ZN(vscale_core_DW01_sub_7n163) );
  INV_X4 vscale_core_DW01_sub_7_U432 ( .A(vscale_core_DW01_sub_7n162), .ZN(vscale_core_DW01_sub_7n160) );
  INV_X4 vscale_core_DW01_sub_7_U433 ( .A(vscale_core_DW01_sub_7n143), .ZN(vscale_core_DW01_sub_7n142) );
  INV_X4 vscale_core_DW01_sub_7_U434 ( .A(vscale_core_DW01_sub_7n136), .ZN(vscale_core_DW01_sub_7n134) );
  INV_X4 vscale_core_DW01_sub_7_U435 ( .A(vscale_core_DW01_sub_7n135), .ZN(vscale_core_DW01_sub_7n133) );
  INV_X4 vscale_core_DW01_sub_7_U436 ( .A(vscale_core_DW01_sub_7n131), .ZN(vscale_core_DW01_sub_7n129) );
  INV_X4 vscale_core_DW01_sub_7_U437 ( .A(vscale_core_DW01_sub_7n130), .ZN(vscale_core_DW01_sub_7n195) );
  INV_X4 vscale_core_DW01_sub_7_U438 ( .A(vscale_core_DW01_sub_7n120), .ZN(vscale_core_DW01_sub_7n119) );
  INV_X4 vscale_core_DW01_sub_7_U439 ( .A(vscale_core_DW01_sub_7n118), .ZN(vscale_core_DW01_sub_7n116) );
  INV_X4 vscale_core_DW01_sub_7_U440 ( .A(vscale_core_DW01_sub_7n117), .ZN(vscale_core_DW01_sub_7n193) );
  INV_X4 vscale_core_DW01_sub_7_U441 ( .A(vscale_core_DW01_sub_7n111), .ZN(vscale_core_DW01_sub_7n109) );
  INV_X4 vscale_core_DW01_sub_7_U442 ( .A(vscale_core_DW01_sub_7n110), .ZN(vscale_core_DW01_sub_7n108) );
  INV_X4 vscale_core_DW01_sub_7_U443 ( .A(vscale_core_DW01_sub_7n106), .ZN(vscale_core_DW01_sub_7n104) );
  INV_X4 vscale_core_DW01_sub_7_U444 ( .A(vscale_core_DW01_sub_7n105), .ZN(vscale_core_DW01_sub_7n191) );
;
  vscale_core_DW01_add_7 pipeline_alu_add_17 

  FA_X1 vscale_core_DW01_add_7_U3 ( .A(pipeline_alu_src_b[30]), .B(n6997), .CI(vscale_core_DW01_add_7n30), .CO(vscale_core_DW01_add_7n29), .S(pipeline_alu_N89) );
  FA_X1 vscale_core_DW01_add_7_U4 ( .A(n6557), .B(pipeline_alu_src_a[29]), .CI(vscale_core_DW01_add_7n31), .CO(vscale_core_DW01_add_7n30), .S(pipeline_alu_N88) );
  FA_X1 vscale_core_DW01_add_7_U5 ( .A(pipeline_alu_src_b[28]), .B(n6565), .CI(vscale_core_DW01_add_7n32), .CO(vscale_core_DW01_add_7n31), .S(pipeline_alu_N87) );
  FA_X1 vscale_core_DW01_add_7_U6 ( .A(pipeline_alu_src_b[27]), .B(n6603), .CI(vscale_core_DW01_add_7n33), .CO(vscale_core_DW01_add_7n32), .S(pipeline_alu_N86) );
  XOR2_X2 vscale_core_DW01_add_7_U7 ( .A(vscale_core_DW01_add_7n2), .B(vscale_core_DW01_add_7n36), .Z(pipeline_alu_N85) );
  NAND2_X2 vscale_core_DW01_add_7_U9 ( .A1(vscale_core_DW01_add_7n174), .A2(vscale_core_DW01_add_7n35), .ZN(vscale_core_DW01_add_7n2) );
  XNOR2_X2 vscale_core_DW01_add_7_U13 ( .A(vscale_core_DW01_add_7n41), .B(vscale_core_DW01_add_7n3), .ZN(pipeline_alu_N84) );
  NAND2_X2 vscale_core_DW01_add_7_U17 ( .A1(vscale_core_DW01_add_7n308), .A2(vscale_core_DW01_add_7n40), .ZN(vscale_core_DW01_add_7n3) );
  NAND2_X2 vscale_core_DW01_add_7_U20 ( .A1(pipeline_alu_src_b[25]), .A2(n6608), .ZN(vscale_core_DW01_add_7n40) );
  XOR2_X2 vscale_core_DW01_add_7_U21 ( .A(vscale_core_DW01_add_7n4), .B(vscale_core_DW01_add_7n44), .Z(pipeline_alu_N83) );
  NAND2_X2 vscale_core_DW01_add_7_U23 ( .A1(vscale_core_DW01_add_7n176), .A2(vscale_core_DW01_add_7n43), .ZN(vscale_core_DW01_add_7n4) );
  NAND2_X2 vscale_core_DW01_add_7_U26 ( .A1(pipeline_alu_src_b[24]), .A2(pipeline_alu_src_a[24]), .ZN(vscale_core_DW01_add_7n43) );
  XNOR2_X2 vscale_core_DW01_add_7_U27 ( .A(vscale_core_DW01_add_7n49), .B(vscale_core_DW01_add_7n5), .ZN(pipeline_alu_N82) );
  NAND2_X2 vscale_core_DW01_add_7_U31 ( .A1(vscale_core_DW01_add_7n307), .A2(vscale_core_DW01_add_7n48), .ZN(vscale_core_DW01_add_7n5) );
  NAND2_X2 vscale_core_DW01_add_7_U34 ( .A1(pipeline_alu_src_b[23]), .A2(n6980), .ZN(vscale_core_DW01_add_7n48) );
  XOR2_X2 vscale_core_DW01_add_7_U35 ( .A(vscale_core_DW01_add_7n6), .B(vscale_core_DW01_add_7n52), .Z(pipeline_alu_N81) );
  NAND2_X2 vscale_core_DW01_add_7_U37 ( .A1(vscale_core_DW01_add_7n178), .A2(vscale_core_DW01_add_7n51), .ZN(vscale_core_DW01_add_7n6) );
  XNOR2_X2 vscale_core_DW01_add_7_U41 ( .A(vscale_core_DW01_add_7n57), .B(vscale_core_DW01_add_7n7), .ZN(pipeline_alu_N80) );
  NAND2_X2 vscale_core_DW01_add_7_U45 ( .A1(vscale_core_DW01_add_7n306), .A2(vscale_core_DW01_add_7n56), .ZN(vscale_core_DW01_add_7n7) );
  XOR2_X2 vscale_core_DW01_add_7_U49 ( .A(vscale_core_DW01_add_7n8), .B(vscale_core_DW01_add_7n64), .Z(pipeline_alu_N79) );
  NAND2_X2 vscale_core_DW01_add_7_U51 ( .A1(vscale_core_DW01_add_7n65), .A2(vscale_core_DW01_add_7n304), .ZN(vscale_core_DW01_add_7n58) );
  NAND2_X2 vscale_core_DW01_add_7_U58 ( .A1(pipeline_alu_src_b[20]), .A2(pipeline_alu_src_a[20]), .ZN(vscale_core_DW01_add_7n63) );
  XOR2_X2 vscale_core_DW01_add_7_U59 ( .A(vscale_core_DW01_add_7n9), .B(vscale_core_DW01_add_7n69), .Z(pipeline_alu_N78) );
  NAND2_X2 vscale_core_DW01_add_7_U63 ( .A1(vscale_core_DW01_add_7n181), .A2(vscale_core_DW01_add_7n68), .ZN(vscale_core_DW01_add_7n9) );
  NAND2_X2 vscale_core_DW01_add_7_U66 ( .A1(pipeline_alu_src_b[19]), .A2(pipeline_alu_src_a[19]), .ZN(vscale_core_DW01_add_7n68) );
  XOR2_X2 vscale_core_DW01_add_7_U67 ( .A(vscale_core_DW01_add_7n10), .B(vscale_core_DW01_add_7n78), .Z(pipeline_alu_N77) );
  NAND2_X2 vscale_core_DW01_add_7_U71 ( .A1(vscale_core_DW01_add_7n79), .A2(vscale_core_DW01_add_7n305), .ZN(vscale_core_DW01_add_7n72) );
  NAND2_X2 vscale_core_DW01_add_7_U78 ( .A1(pipeline_alu_src_b[18]), .A2(pipeline_alu_src_a[18]), .ZN(vscale_core_DW01_add_7n77) );
  XOR2_X2 vscale_core_DW01_add_7_U79 ( .A(vscale_core_DW01_add_7n11), .B(vscale_core_DW01_add_7n83), .Z(pipeline_alu_N76) );
  NAND2_X2 vscale_core_DW01_add_7_U83 ( .A1(vscale_core_DW01_add_7n183), .A2(vscale_core_DW01_add_7n82), .ZN(vscale_core_DW01_add_7n11) );
  XNOR2_X2 vscale_core_DW01_add_7_U87 ( .A(vscale_core_DW01_add_7n88), .B(vscale_core_DW01_add_7n12), .ZN(pipeline_alu_N75) );
  NAND2_X2 vscale_core_DW01_add_7_U91 ( .A1(vscale_core_DW01_add_7n84), .A2(vscale_core_DW01_add_7n87), .ZN(vscale_core_DW01_add_7n12) );
  XOR2_X2 vscale_core_DW01_add_7_U95 ( .A(vscale_core_DW01_add_7n13), .B(vscale_core_DW01_add_7n98), .Z(pipeline_alu_N74) );
  NAND2_X2 vscale_core_DW01_add_7_U100 ( .A1(vscale_core_DW01_add_7n106), .A2(vscale_core_DW01_add_7n94), .ZN(vscale_core_DW01_add_7n92) );
  NAND2_X2 vscale_core_DW01_add_7_U104 ( .A1(vscale_core_DW01_add_7n185), .A2(vscale_core_DW01_add_7n97), .ZN(vscale_core_DW01_add_7n13) );
  XNOR2_X2 vscale_core_DW01_add_7_U108 ( .A(vscale_core_DW01_add_7n103), .B(vscale_core_DW01_add_7n14), .ZN(pipeline_alu_N73) );
  NAND2_X2 vscale_core_DW01_add_7_U112 ( .A1(vscale_core_DW01_add_7n99), .A2(vscale_core_DW01_add_7n102), .ZN(vscale_core_DW01_add_7n14) );
  XOR2_X2 vscale_core_DW01_add_7_U116 ( .A(vscale_core_DW01_add_7n15), .B(vscale_core_DW01_add_7n110), .Z(pipeline_alu_N72) );
  NAND2_X2 vscale_core_DW01_add_7_U122 ( .A1(vscale_core_DW01_add_7n187), .A2(vscale_core_DW01_add_7n109), .ZN(vscale_core_DW01_add_7n15) );
  XOR2_X2 vscale_core_DW01_add_7_U126 ( .A(vscale_core_DW01_add_7n16), .B(vscale_core_DW01_add_7n115), .Z(pipeline_alu_N71) );
  NAND2_X2 vscale_core_DW01_add_7_U130 ( .A1(vscale_core_DW01_add_7n188), .A2(vscale_core_DW01_add_7n114), .ZN(vscale_core_DW01_add_7n16) );
  XOR2_X2 vscale_core_DW01_add_7_U134 ( .A(vscale_core_DW01_add_7n17), .B(vscale_core_DW01_add_7n123), .Z(pipeline_alu_N70) );
  NAND2_X2 vscale_core_DW01_add_7_U137 ( .A1(vscale_core_DW01_add_7n131), .A2(vscale_core_DW01_add_7n119), .ZN(vscale_core_DW01_add_7n117) );
  NAND2_X2 vscale_core_DW01_add_7_U141 ( .A1(vscale_core_DW01_add_7n189), .A2(vscale_core_DW01_add_7n122), .ZN(vscale_core_DW01_add_7n17) );
  XNOR2_X2 vscale_core_DW01_add_7_U145 ( .A(vscale_core_DW01_add_7n128), .B(vscale_core_DW01_add_7n18), .ZN(pipeline_alu_N69) );
  NAND2_X2 vscale_core_DW01_add_7_U149 ( .A1(vscale_core_DW01_add_7n190), .A2(vscale_core_DW01_add_7n127), .ZN(vscale_core_DW01_add_7n18) );
  XNOR2_X2 vscale_core_DW01_add_7_U153 ( .A(vscale_core_DW01_add_7n135), .B(vscale_core_DW01_add_7n19), .ZN(pipeline_alu_N68) );
  NAND2_X2 vscale_core_DW01_add_7_U159 ( .A1(vscale_core_DW01_add_7n191), .A2(vscale_core_DW01_add_7n134), .ZN(vscale_core_DW01_add_7n19) );
  NAND2_X2 vscale_core_DW01_add_7_U162 ( .A1(n6973), .A2(pipeline_alu_src_b[9]), .ZN(vscale_core_DW01_add_7n134) );
  XOR2_X2 vscale_core_DW01_add_7_U163 ( .A(vscale_core_DW01_add_7n20), .B(vscale_core_DW01_add_7n138), .Z(pipeline_alu_N67) );
  NAND2_X2 vscale_core_DW01_add_7_U165 ( .A1(vscale_core_DW01_add_7n192), .A2(vscale_core_DW01_add_7n137), .ZN(vscale_core_DW01_add_7n20) );
  XNOR2_X2 vscale_core_DW01_add_7_U169 ( .A(vscale_core_DW01_add_7n146), .B(vscale_core_DW01_add_7n21), .ZN(pipeline_alu_N66) );
  NAND2_X2 vscale_core_DW01_add_7_U172 ( .A1(vscale_core_DW01_add_7n150), .A2(vscale_core_DW01_add_7n142), .ZN(vscale_core_DW01_add_7n140) );
  NAND2_X2 vscale_core_DW01_add_7_U176 ( .A1(vscale_core_DW01_add_7n193), .A2(vscale_core_DW01_add_7n145), .ZN(vscale_core_DW01_add_7n21) );
  XOR2_X2 vscale_core_DW01_add_7_U180 ( .A(vscale_core_DW01_add_7n22), .B(vscale_core_DW01_add_7n149), .Z(pipeline_alu_N65) );
  NAND2_X2 vscale_core_DW01_add_7_U182 ( .A1(vscale_core_DW01_add_7n194), .A2(vscale_core_DW01_add_7n148), .ZN(vscale_core_DW01_add_7n22) );
  XOR2_X2 vscale_core_DW01_add_7_U186 ( .A(vscale_core_DW01_add_7n23), .B(vscale_core_DW01_add_7n154), .Z(pipeline_alu_N64) );
  NAND2_X2 vscale_core_DW01_add_7_U190 ( .A1(vscale_core_DW01_add_7n195), .A2(vscale_core_DW01_add_7n153), .ZN(vscale_core_DW01_add_7n23) );
  XNOR2_X2 vscale_core_DW01_add_7_U194 ( .A(vscale_core_DW01_add_7n159), .B(vscale_core_DW01_add_7n24), .ZN(pipeline_alu_N63) );
  XNOR2_X2 vscale_core_DW01_add_7_U202 ( .A(vscale_core_DW01_add_7n165), .B(vscale_core_DW01_add_7n25), .ZN(pipeline_alu_N62) );
  NAND2_X2 vscale_core_DW01_add_7_U207 ( .A1(vscale_core_DW01_add_7n197), .A2(vscale_core_DW01_add_7n164), .ZN(vscale_core_DW01_add_7n25) );
  XOR2_X2 vscale_core_DW01_add_7_U211 ( .A(vscale_core_DW01_add_7n26), .B(vscale_core_DW01_add_7n168), .Z(pipeline_alu_N61) );
  NAND2_X2 vscale_core_DW01_add_7_U213 ( .A1(vscale_core_DW01_add_7n198), .A2(vscale_core_DW01_add_7n167), .ZN(vscale_core_DW01_add_7n26) );
  XOR2_X2 vscale_core_DW01_add_7_U217 ( .A(vscale_core_DW01_add_7n173), .B(vscale_core_DW01_add_7n27), .Z(pipeline_alu_N60) );
  NAND2_X2 vscale_core_DW01_add_7_U220 ( .A1(vscale_core_DW01_add_7n199), .A2(vscale_core_DW01_add_7n171), .ZN(vscale_core_DW01_add_7n27) );
  NAND2_X1 vscale_core_DW01_add_7_U232 ( .A1(pipeline_alu_src_b[13]), .A2(n6566), .ZN(vscale_core_DW01_add_7n109) );
  NAND2_X1 vscale_core_DW01_add_7_U233 ( .A1(pipeline_alu_src_b[26]), .A2(n6560), .ZN(vscale_core_DW01_add_7n35) );
  AOI21_X2 vscale_core_DW01_add_7_U234 ( .B1(vscale_core_DW01_add_7n57), .B2(vscale_core_DW01_add_7n306), .A(vscale_core_DW01_add_7n54), .ZN(vscale_core_DW01_add_7n52) );
  XOR2_X1 vscale_core_DW01_add_7_U235 ( .A(n13159), .B(n7006), .Z(vscale_core_DW01_add_7n1) );
  NAND2_X1 vscale_core_DW01_add_7_U236 ( .A1(pipeline_alu_src_b[22]), .A2(n6626), .ZN(vscale_core_DW01_add_7n51) );
  AOI21_X2 vscale_core_DW01_add_7_U237 ( .B1(vscale_core_DW01_add_7n49), .B2(vscale_core_DW01_add_7n307), .A(vscale_core_DW01_add_7n46), .ZN(vscale_core_DW01_add_7n44) );
  AND2_X4 vscale_core_DW01_add_7_U238 ( .A1(vscale_core_DW01_add_7n309), .A2(vscale_core_DW01_add_7n173), .ZN(pipeline_alu_N59) );
  NAND2_X1 vscale_core_DW01_add_7_U239 ( .A1(pipeline_alu_src_b[21]), .A2(pipeline_alu_src_a[21]), .ZN(vscale_core_DW01_add_7n56) );
  NAND2_X1 vscale_core_DW01_add_7_U240 ( .A1(n9398), .A2(pipeline_alu_src_a[2]), .ZN(vscale_core_DW01_add_7n167) );
  NAND2_X1 vscale_core_DW01_add_7_U241 ( .A1(n6618), .A2(pipeline_alu_src_a[0]), .ZN(vscale_core_DW01_add_7n173) );
  NAND2_X1 vscale_core_DW01_add_7_U242 ( .A1(n6620), .A2(pipeline_alu_src_b[5]), .ZN(vscale_core_DW01_add_7n153) );
  NAND2_X1 vscale_core_DW01_add_7_U243 ( .A1(n6614), .A2(pipeline_alu_src_b[11]), .ZN(vscale_core_DW01_add_7n122) );
  NAND2_X1 vscale_core_DW01_add_7_U244 ( .A1(pipeline_alu_src_b[17]), .A2(pipeline_alu_src_a[17]), .ZN(vscale_core_DW01_add_7n82) );
  NAND2_X1 vscale_core_DW01_add_7_U245 ( .A1(n6600), .A2(pipeline_alu_src_a[4]), .ZN(vscale_core_DW01_add_7n158) );
  NAND2_X1 vscale_core_DW01_add_7_U246 ( .A1(vscale_core_DW01_add_7n196), .A2(vscale_core_DW01_add_7n158), .ZN(vscale_core_DW01_add_7n24) );
  INV_X1 vscale_core_DW01_add_7_U247 ( .A(vscale_core_DW01_add_7n158), .ZN(vscale_core_DW01_add_7n156) );
  NOR2_X2 vscale_core_DW01_add_7_U248 ( .A1(vscale_core_DW01_add_7n113), .A2(vscale_core_DW01_add_7n108), .ZN(vscale_core_DW01_add_7n106) );
  NOR2_X2 vscale_core_DW01_add_7_U249 ( .A1(vscale_core_DW01_add_7n72), .A2(vscale_core_DW01_add_7n67), .ZN(vscale_core_DW01_add_7n65) );
  AOI21_X4 vscale_core_DW01_add_7_U250 ( .B1(vscale_core_DW01_add_7n139), .B2(vscale_core_DW01_add_7n90), .A(vscale_core_DW01_add_7n91), .ZN(vscale_core_DW01_add_7n89) );
  NOR2_X1 vscale_core_DW01_add_7_U251 ( .A1(vscale_core_DW01_add_7n92), .A2(vscale_core_DW01_add_7n117), .ZN(vscale_core_DW01_add_7n90) );
  NOR2_X1 vscale_core_DW01_add_7_U252 ( .A1(vscale_core_DW01_add_7n147), .A2(vscale_core_DW01_add_7n144), .ZN(vscale_core_DW01_add_7n142) );
  OAI21_X1 vscale_core_DW01_add_7_U253 ( .B1(vscale_core_DW01_add_7n133), .B2(vscale_core_DW01_add_7n137), .A(vscale_core_DW01_add_7n134), .ZN(vscale_core_DW01_add_7n132) );
  OAI21_X1 vscale_core_DW01_add_7_U254 ( .B1(vscale_core_DW01_add_7n170), .B2(vscale_core_DW01_add_7n173), .A(vscale_core_DW01_add_7n171), .ZN(vscale_core_DW01_add_7n169) );
  OAI21_X1 vscale_core_DW01_add_7_U255 ( .B1(vscale_core_DW01_add_7n81), .B2(vscale_core_DW01_add_7n87), .A(vscale_core_DW01_add_7n82), .ZN(vscale_core_DW01_add_7n80) );
  OAI21_X1 vscale_core_DW01_add_7_U256 ( .B1(vscale_core_DW01_add_7n152), .B2(vscale_core_DW01_add_7n158), .A(vscale_core_DW01_add_7n153), .ZN(vscale_core_DW01_add_7n151) );
  NOR2_X1 vscale_core_DW01_add_7_U257 ( .A1(vscale_core_DW01_add_7n136), .A2(vscale_core_DW01_add_7n133), .ZN(vscale_core_DW01_add_7n131) );
  NOR2_X1 vscale_core_DW01_add_7_U258 ( .A1(vscale_core_DW01_add_7n81), .A2(vscale_core_DW01_add_7n86), .ZN(vscale_core_DW01_add_7n79) );
  NOR2_X1 vscale_core_DW01_add_7_U259 ( .A1(vscale_core_DW01_add_7n157), .A2(vscale_core_DW01_add_7n152), .ZN(vscale_core_DW01_add_7n150) );
  INV_X1 vscale_core_DW01_add_7_U260 ( .A(vscale_core_DW01_add_7n96), .ZN(vscale_core_DW01_add_7n185) );
  AOI21_X1 vscale_core_DW01_add_7_U261 ( .B1(vscale_core_DW01_add_7n88), .B2(vscale_core_DW01_add_7n65), .A(vscale_core_DW01_add_7n66), .ZN(vscale_core_DW01_add_7n64) );
  NAND2_X1 vscale_core_DW01_add_7_U262 ( .A1(vscale_core_DW01_add_7n304), .A2(vscale_core_DW01_add_7n63), .ZN(vscale_core_DW01_add_7n8) );
  INV_X1 vscale_core_DW01_add_7_U263 ( .A(vscale_core_DW01_add_7n152), .ZN(vscale_core_DW01_add_7n195) );
  INV_X1 vscale_core_DW01_add_7_U264 ( .A(vscale_core_DW01_add_7n108), .ZN(vscale_core_DW01_add_7n187) );
  INV_X1 vscale_core_DW01_add_7_U265 ( .A(vscale_core_DW01_add_7n81), .ZN(vscale_core_DW01_add_7n183) );
  AOI21_X1 vscale_core_DW01_add_7_U266 ( .B1(vscale_core_DW01_add_7n88), .B2(vscale_core_DW01_add_7n79), .A(vscale_core_DW01_add_7n80), .ZN(vscale_core_DW01_add_7n78) );
  NAND2_X1 vscale_core_DW01_add_7_U267 ( .A1(vscale_core_DW01_add_7n305), .A2(vscale_core_DW01_add_7n77), .ZN(vscale_core_DW01_add_7n10) );
  INV_X1 vscale_core_DW01_add_7_U268 ( .A(vscale_core_DW01_add_7n67), .ZN(vscale_core_DW01_add_7n181) );
  OAI21_X1 vscale_core_DW01_add_7_U269 ( .B1(vscale_core_DW01_add_7n149), .B2(vscale_core_DW01_add_7n147), .A(vscale_core_DW01_add_7n148), .ZN(vscale_core_DW01_add_7n146) );
  INV_X1 vscale_core_DW01_add_7_U270 ( .A(vscale_core_DW01_add_7n144), .ZN(vscale_core_DW01_add_7n193) );
  INV_X1 vscale_core_DW01_add_7_U271 ( .A(vscale_core_DW01_add_7n133), .ZN(vscale_core_DW01_add_7n191) );
  INV_X1 vscale_core_DW01_add_7_U272 ( .A(vscale_core_DW01_add_7n163), .ZN(vscale_core_DW01_add_7n197) );
  INV_X1 vscale_core_DW01_add_7_U273 ( .A(vscale_core_DW01_add_7n86), .ZN(vscale_core_DW01_add_7n84) );
  INV_X1 vscale_core_DW01_add_7_U274 ( .A(vscale_core_DW01_add_7n121), .ZN(vscale_core_DW01_add_7n189) );
  NOR2_X1 vscale_core_DW01_add_7_U275 ( .A1(vscale_core_DW01_add_7n126), .A2(vscale_core_DW01_add_7n121), .ZN(vscale_core_DW01_add_7n119) );
  XOR2_X1 vscale_core_DW01_add_7_U276 ( .A(vscale_core_DW01_add_7n1), .B(vscale_core_DW01_add_7n29), .Z(pipeline_alu_N90) );
  OAI21_X2 vscale_core_DW01_add_7_U277 ( .B1(vscale_core_DW01_add_7n118), .B2(vscale_core_DW01_add_7n92), .A(vscale_core_DW01_add_7n93), .ZN(vscale_core_DW01_add_7n91) );
  AOI21_X2 vscale_core_DW01_add_7_U278 ( .B1(vscale_core_DW01_add_7n159), .B2(vscale_core_DW01_add_7n150), .A(vscale_core_DW01_add_7n151), .ZN(vscale_core_DW01_add_7n149) );
  OAI21_X1 vscale_core_DW01_add_7_U279 ( .B1(vscale_core_DW01_add_7n138), .B2(vscale_core_DW01_add_7n117), .A(vscale_core_DW01_add_7n118), .ZN(vscale_core_DW01_add_7n116) );
  OAI21_X2 vscale_core_DW01_add_7_U280 ( .B1(vscale_core_DW01_add_7n138), .B2(vscale_core_DW01_add_7n129), .A(vscale_core_DW01_add_7n130), .ZN(vscale_core_DW01_add_7n128) );
  OAI21_X2 vscale_core_DW01_add_7_U281 ( .B1(vscale_core_DW01_add_7n115), .B2(vscale_core_DW01_add_7n104), .A(vscale_core_DW01_add_7n105), .ZN(vscale_core_DW01_add_7n103) );
  AOI21_X2 vscale_core_DW01_add_7_U282 ( .B1(vscale_core_DW01_add_7n41), .B2(vscale_core_DW01_add_7n308), .A(vscale_core_DW01_add_7n38), .ZN(vscale_core_DW01_add_7n36) );
  AOI21_X2 vscale_core_DW01_add_7_U283 ( .B1(vscale_core_DW01_add_7n119), .B2(vscale_core_DW01_add_7n132), .A(vscale_core_DW01_add_7n120), .ZN(vscale_core_DW01_add_7n118) );
  OAI21_X1 vscale_core_DW01_add_7_U284 ( .B1(vscale_core_DW01_add_7n121), .B2(vscale_core_DW01_add_7n127), .A(vscale_core_DW01_add_7n122), .ZN(vscale_core_DW01_add_7n120) );
  AOI21_X2 vscale_core_DW01_add_7_U285 ( .B1(vscale_core_DW01_add_7n80), .B2(vscale_core_DW01_add_7n305), .A(vscale_core_DW01_add_7n75), .ZN(vscale_core_DW01_add_7n73) );
  AOI21_X2 vscale_core_DW01_add_7_U286 ( .B1(vscale_core_DW01_add_7n161), .B2(vscale_core_DW01_add_7n169), .A(vscale_core_DW01_add_7n162), .ZN(vscale_core_DW01_add_7n160) );
  NOR2_X2 vscale_core_DW01_add_7_U287 ( .A1(vscale_core_DW01_add_7n166), .A2(vscale_core_DW01_add_7n163), .ZN(vscale_core_DW01_add_7n161) );
  OAI21_X2 vscale_core_DW01_add_7_U288 ( .B1(vscale_core_DW01_add_7n163), .B2(vscale_core_DW01_add_7n167), .A(vscale_core_DW01_add_7n164), .ZN(vscale_core_DW01_add_7n162) );
  OAI21_X2 vscale_core_DW01_add_7_U289 ( .B1(vscale_core_DW01_add_7n73), .B2(vscale_core_DW01_add_7n67), .A(vscale_core_DW01_add_7n68), .ZN(vscale_core_DW01_add_7n66) );
  OAI21_X2 vscale_core_DW01_add_7_U290 ( .B1(vscale_core_DW01_add_7n160), .B2(vscale_core_DW01_add_7n140), .A(vscale_core_DW01_add_7n141), .ZN(vscale_core_DW01_add_7n139) );
  AOI21_X2 vscale_core_DW01_add_7_U291 ( .B1(vscale_core_DW01_add_7n151), .B2(vscale_core_DW01_add_7n142), .A(vscale_core_DW01_add_7n143), .ZN(vscale_core_DW01_add_7n141) );
  OAI21_X2 vscale_core_DW01_add_7_U292 ( .B1(vscale_core_DW01_add_7n52), .B2(vscale_core_DW01_add_7n50), .A(vscale_core_DW01_add_7n51), .ZN(vscale_core_DW01_add_7n49) );
  OAI21_X2 vscale_core_DW01_add_7_U293 ( .B1(vscale_core_DW01_add_7n44), .B2(vscale_core_DW01_add_7n42), .A(vscale_core_DW01_add_7n43), .ZN(vscale_core_DW01_add_7n41) );
  OAI21_X2 vscale_core_DW01_add_7_U294 ( .B1(vscale_core_DW01_add_7n89), .B2(vscale_core_DW01_add_7n58), .A(vscale_core_DW01_add_7n59), .ZN(vscale_core_DW01_add_7n57) );
  AOI21_X2 vscale_core_DW01_add_7_U295 ( .B1(vscale_core_DW01_add_7n66), .B2(vscale_core_DW01_add_7n304), .A(vscale_core_DW01_add_7n61), .ZN(vscale_core_DW01_add_7n59) );
  OAI21_X2 vscale_core_DW01_add_7_U296 ( .B1(vscale_core_DW01_add_7n108), .B2(vscale_core_DW01_add_7n114), .A(vscale_core_DW01_add_7n109), .ZN(vscale_core_DW01_add_7n107) );
  AOI21_X2 vscale_core_DW01_add_7_U297 ( .B1(vscale_core_DW01_add_7n94), .B2(vscale_core_DW01_add_7n107), .A(vscale_core_DW01_add_7n95), .ZN(vscale_core_DW01_add_7n93) );
  OAI21_X1 vscale_core_DW01_add_7_U298 ( .B1(vscale_core_DW01_add_7n96), .B2(vscale_core_DW01_add_7n102), .A(vscale_core_DW01_add_7n97), .ZN(vscale_core_DW01_add_7n95) );
  OAI21_X1 vscale_core_DW01_add_7_U299 ( .B1(vscale_core_DW01_add_7n144), .B2(vscale_core_DW01_add_7n148), .A(vscale_core_DW01_add_7n145), .ZN(vscale_core_DW01_add_7n143) );
  NOR2_X1 vscale_core_DW01_add_7_U300 ( .A1(vscale_core_DW01_add_7n101), .A2(vscale_core_DW01_add_7n96), .ZN(vscale_core_DW01_add_7n94) );
  AOI21_X2 vscale_core_DW01_add_7_U301 ( .B1(vscale_core_DW01_add_7n159), .B2(vscale_core_DW01_add_7n196), .A(vscale_core_DW01_add_7n156), .ZN(vscale_core_DW01_add_7n154) );
  AOI21_X2 vscale_core_DW01_add_7_U302 ( .B1(vscale_core_DW01_add_7n128), .B2(vscale_core_DW01_add_7n190), .A(vscale_core_DW01_add_7n125), .ZN(vscale_core_DW01_add_7n123) );
  AOI21_X2 vscale_core_DW01_add_7_U303 ( .B1(vscale_core_DW01_add_7n116), .B2(vscale_core_DW01_add_7n188), .A(vscale_core_DW01_add_7n112), .ZN(vscale_core_DW01_add_7n110) );
  AOI21_X2 vscale_core_DW01_add_7_U304 ( .B1(vscale_core_DW01_add_7n103), .B2(vscale_core_DW01_add_7n99), .A(vscale_core_DW01_add_7n100), .ZN(vscale_core_DW01_add_7n98) );
  AOI21_X2 vscale_core_DW01_add_7_U305 ( .B1(vscale_core_DW01_add_7n88), .B2(vscale_core_DW01_add_7n84), .A(vscale_core_DW01_add_7n85), .ZN(vscale_core_DW01_add_7n83) );
  AOI21_X2 vscale_core_DW01_add_7_U306 ( .B1(vscale_core_DW01_add_7n88), .B2(vscale_core_DW01_add_7n70), .A(vscale_core_DW01_add_7n71), .ZN(vscale_core_DW01_add_7n69) );
  OAI21_X1 vscale_core_DW01_add_7_U307 ( .B1(vscale_core_DW01_add_7n138), .B2(vscale_core_DW01_add_7n136), .A(vscale_core_DW01_add_7n137), .ZN(vscale_core_DW01_add_7n135) );
  OAI21_X1 vscale_core_DW01_add_7_U308 ( .B1(vscale_core_DW01_add_7n168), .B2(vscale_core_DW01_add_7n166), .A(vscale_core_DW01_add_7n167), .ZN(vscale_core_DW01_add_7n165) );
  NOR2_X1 vscale_core_DW01_add_7_U309 ( .A1(pipeline_alu_src_b[17]), .A2(pipeline_alu_src_a[17]), .ZN(vscale_core_DW01_add_7n81) );
  NOR2_X1 vscale_core_DW01_add_7_U310 ( .A1(pipeline_alu_src_b[13]), .A2(n6566), .ZN(vscale_core_DW01_add_7n108) );
  NOR2_X1 vscale_core_DW01_add_7_U311 ( .A1(n6620), .A2(pipeline_alu_src_b[5]), .ZN(vscale_core_DW01_add_7n152) );
  NOR2_X1 vscale_core_DW01_add_7_U312 ( .A1(n6973), .A2(pipeline_alu_src_b[9]), .ZN(vscale_core_DW01_add_7n133) );
  NOR2_X1 vscale_core_DW01_add_7_U313 ( .A1(n6614), .A2(pipeline_alu_src_b[11]), .ZN(vscale_core_DW01_add_7n121) );
  OAI21_X2 vscale_core_DW01_add_7_U314 ( .B1(vscale_core_DW01_add_7n36), .B2(vscale_core_DW01_add_7n34), .A(vscale_core_DW01_add_7n35), .ZN(vscale_core_DW01_add_7n33) );
  NOR2_X1 vscale_core_DW01_add_7_U315 ( .A1(pipeline_alu_src_b[19]), .A2(pipeline_alu_src_a[19]), .ZN(vscale_core_DW01_add_7n67) );
  NOR2_X1 vscale_core_DW01_add_7_U316 ( .A1(n9398), .A2(pipeline_alu_src_a[2]), .ZN(vscale_core_DW01_add_7n166) );
  NOR2_X1 vscale_core_DW01_add_7_U317 ( .A1(n6600), .A2(pipeline_alu_src_a[4]), .ZN(vscale_core_DW01_add_7n157) );
  OR2_X1 vscale_core_DW01_add_7_U318 ( .A1(pipeline_alu_src_b[20]), .A2(pipeline_alu_src_a[20]), .ZN(vscale_core_DW01_add_7n304) );
  OR2_X1 vscale_core_DW01_add_7_U319 ( .A1(pipeline_alu_src_b[18]), .A2(pipeline_alu_src_a[18]), .ZN(vscale_core_DW01_add_7n305) );
  OR2_X1 vscale_core_DW01_add_7_U320 ( .A1(pipeline_alu_src_b[21]), .A2(pipeline_alu_src_a[21]), .ZN(vscale_core_DW01_add_7n306) );
  NOR2_X1 vscale_core_DW01_add_7_U321 ( .A1(pipeline_alu_src_b[22]), .A2(n6626), .ZN(vscale_core_DW01_add_7n50) );
  NOR2_X1 vscale_core_DW01_add_7_U322 ( .A1(pipeline_alu_src_b[24]), .A2(pipeline_alu_src_a[24]), .ZN(vscale_core_DW01_add_7n42) );
  NOR2_X1 vscale_core_DW01_add_7_U323 ( .A1(pipeline_alu_src_b[26]), .A2(n6560), .ZN(vscale_core_DW01_add_7n34) );
  OR2_X1 vscale_core_DW01_add_7_U324 ( .A1(pipeline_alu_src_b[23]), .A2(n6980), .ZN(vscale_core_DW01_add_7n307) );
  OR2_X1 vscale_core_DW01_add_7_U325 ( .A1(pipeline_alu_src_b[25]), .A2(n6608), .ZN(vscale_core_DW01_add_7n308) );
  OR2_X1 vscale_core_DW01_add_7_U326 ( .A1(n6618), .A2(pipeline_alu_src_a[0]), .ZN(vscale_core_DW01_add_7n309) );
  NOR2_X1 vscale_core_DW01_add_7_U327 ( .A1(n6929), .A2(n6634), .ZN(vscale_core_DW01_add_7n163) );
  NOR2_X1 vscale_core_DW01_add_7_U328 ( .A1(n6571), .A2(pipeline_alu_src_b[10]), .ZN(vscale_core_DW01_add_7n126) );
  NAND2_X1 vscale_core_DW01_add_7_U329 ( .A1(n6571), .A2(pipeline_alu_src_b[10]), .ZN(vscale_core_DW01_add_7n127) );
  NAND2_X1 vscale_core_DW01_add_7_U330 ( .A1(pipeline_alu_src_b[14]), .A2(pipeline_alu_src_a[14]), .ZN(vscale_core_DW01_add_7n102) );
  NOR2_X1 vscale_core_DW01_add_7_U331 ( .A1(pipeline_alu_src_b[14]), .A2(pipeline_alu_src_a[14]), .ZN(vscale_core_DW01_add_7n101) );
  NOR2_X1 vscale_core_DW01_add_7_U332 ( .A1(n6976), .A2(pipeline_alu_src_a[1]), .ZN(vscale_core_DW01_add_7n170) );
  NAND2_X1 vscale_core_DW01_add_7_U333 ( .A1(n6976), .A2(pipeline_alu_src_a[1]), .ZN(vscale_core_DW01_add_7n171) );
  NAND2_X1 vscale_core_DW01_add_7_U334 ( .A1(n6611), .A2(pipeline_alu_src_b[7]), .ZN(vscale_core_DW01_add_7n145) );
  NOR2_X1 vscale_core_DW01_add_7_U335 ( .A1(n6611), .A2(pipeline_alu_src_b[7]), .ZN(vscale_core_DW01_add_7n144) );
  NOR2_X1 vscale_core_DW01_add_7_U336 ( .A1(pipeline_alu_src_b[12]), .A2(pipeline_alu_src_a[12]), .ZN(vscale_core_DW01_add_7n113) );
  NAND2_X1 vscale_core_DW01_add_7_U337 ( .A1(pipeline_alu_src_b[12]), .A2(pipeline_alu_src_a[12]), .ZN(vscale_core_DW01_add_7n114) );
  NAND2_X1 vscale_core_DW01_add_7_U338 ( .A1(pipeline_alu_src_b[15]), .A2(n6597), .ZN(vscale_core_DW01_add_7n97) );
  NOR2_X1 vscale_core_DW01_add_7_U339 ( .A1(pipeline_alu_src_b[15]), .A2(n6597), .ZN(vscale_core_DW01_add_7n96) );
  NOR2_X1 vscale_core_DW01_add_7_U340 ( .A1(pipeline_alu_src_b[16]), .A2(pipeline_alu_src_a[16]), .ZN(vscale_core_DW01_add_7n86) );
  NAND2_X1 vscale_core_DW01_add_7_U341 ( .A1(pipeline_alu_src_b[16]), .A2(pipeline_alu_src_a[16]), .ZN(vscale_core_DW01_add_7n87) );
  NOR2_X1 vscale_core_DW01_add_7_U342 ( .A1(n6606), .A2(pipeline_alu_src_b[6]), .ZN(vscale_core_DW01_add_7n147) );
  NAND2_X1 vscale_core_DW01_add_7_U343 ( .A1(n6606), .A2(pipeline_alu_src_b[6]), .ZN(vscale_core_DW01_add_7n148) );
  NOR2_X1 vscale_core_DW01_add_7_U344 ( .A1(n9335), .A2(pipeline_alu_src_b[8]), .ZN(vscale_core_DW01_add_7n136) );
  NAND2_X1 vscale_core_DW01_add_7_U345 ( .A1(n9335), .A2(pipeline_alu_src_b[8]), .ZN(vscale_core_DW01_add_7n137) );
  NAND2_X1 vscale_core_DW01_add_7_U346 ( .A1(n6929), .A2(n6634), .ZN(vscale_core_DW01_add_7n164) );
  INV_X4 vscale_core_DW01_add_7_U347 ( .A(vscale_core_DW01_add_7n89), .ZN(vscale_core_DW01_add_7n88) );
  INV_X4 vscale_core_DW01_add_7_U348 ( .A(vscale_core_DW01_add_7n87), .ZN(vscale_core_DW01_add_7n85) );
  INV_X4 vscale_core_DW01_add_7_U349 ( .A(vscale_core_DW01_add_7n77), .ZN(vscale_core_DW01_add_7n75) );
  INV_X4 vscale_core_DW01_add_7_U350 ( .A(vscale_core_DW01_add_7n73), .ZN(vscale_core_DW01_add_7n71) );
  INV_X4 vscale_core_DW01_add_7_U351 ( .A(vscale_core_DW01_add_7n72), .ZN(vscale_core_DW01_add_7n70) );
  INV_X4 vscale_core_DW01_add_7_U352 ( .A(vscale_core_DW01_add_7n63), .ZN(vscale_core_DW01_add_7n61) );
  INV_X4 vscale_core_DW01_add_7_U353 ( .A(vscale_core_DW01_add_7n56), .ZN(vscale_core_DW01_add_7n54) );
  INV_X4 vscale_core_DW01_add_7_U354 ( .A(vscale_core_DW01_add_7n48), .ZN(vscale_core_DW01_add_7n46) );
  INV_X4 vscale_core_DW01_add_7_U355 ( .A(vscale_core_DW01_add_7n40), .ZN(vscale_core_DW01_add_7n38) );
  INV_X4 vscale_core_DW01_add_7_U356 ( .A(vscale_core_DW01_add_7n170), .ZN(vscale_core_DW01_add_7n199) );
  INV_X4 vscale_core_DW01_add_7_U357 ( .A(vscale_core_DW01_add_7n166), .ZN(vscale_core_DW01_add_7n198) );
  INV_X4 vscale_core_DW01_add_7_U358 ( .A(vscale_core_DW01_add_7n147), .ZN(vscale_core_DW01_add_7n194) );
  INV_X4 vscale_core_DW01_add_7_U359 ( .A(vscale_core_DW01_add_7n136), .ZN(vscale_core_DW01_add_7n192) );
  INV_X4 vscale_core_DW01_add_7_U360 ( .A(vscale_core_DW01_add_7n101), .ZN(vscale_core_DW01_add_7n99) );
  INV_X4 vscale_core_DW01_add_7_U361 ( .A(vscale_core_DW01_add_7n50), .ZN(vscale_core_DW01_add_7n178) );
  INV_X4 vscale_core_DW01_add_7_U362 ( .A(vscale_core_DW01_add_7n42), .ZN(vscale_core_DW01_add_7n176) );
  INV_X4 vscale_core_DW01_add_7_U363 ( .A(vscale_core_DW01_add_7n34), .ZN(vscale_core_DW01_add_7n174) );
  INV_X4 vscale_core_DW01_add_7_U364 ( .A(vscale_core_DW01_add_7n169), .ZN(vscale_core_DW01_add_7n168) );
  INV_X4 vscale_core_DW01_add_7_U365 ( .A(vscale_core_DW01_add_7n160), .ZN(vscale_core_DW01_add_7n159) );
  INV_X4 vscale_core_DW01_add_7_U366 ( .A(vscale_core_DW01_add_7n157), .ZN(vscale_core_DW01_add_7n196) );
  INV_X4 vscale_core_DW01_add_7_U367 ( .A(vscale_core_DW01_add_7n139), .ZN(vscale_core_DW01_add_7n138) );
  INV_X4 vscale_core_DW01_add_7_U368 ( .A(vscale_core_DW01_add_7n132), .ZN(vscale_core_DW01_add_7n130) );
  INV_X4 vscale_core_DW01_add_7_U369 ( .A(vscale_core_DW01_add_7n131), .ZN(vscale_core_DW01_add_7n129) );
  INV_X4 vscale_core_DW01_add_7_U370 ( .A(vscale_core_DW01_add_7n127), .ZN(vscale_core_DW01_add_7n125) );
  INV_X4 vscale_core_DW01_add_7_U371 ( .A(vscale_core_DW01_add_7n126), .ZN(vscale_core_DW01_add_7n190) );
  INV_X4 vscale_core_DW01_add_7_U372 ( .A(vscale_core_DW01_add_7n116), .ZN(vscale_core_DW01_add_7n115) );
  INV_X4 vscale_core_DW01_add_7_U373 ( .A(vscale_core_DW01_add_7n114), .ZN(vscale_core_DW01_add_7n112) );
  INV_X4 vscale_core_DW01_add_7_U374 ( .A(vscale_core_DW01_add_7n113), .ZN(vscale_core_DW01_add_7n188) );
  INV_X4 vscale_core_DW01_add_7_U375 ( .A(vscale_core_DW01_add_7n107), .ZN(vscale_core_DW01_add_7n105) );
  INV_X4 vscale_core_DW01_add_7_U376 ( .A(vscale_core_DW01_add_7n106), .ZN(vscale_core_DW01_add_7n104) );
  INV_X4 vscale_core_DW01_add_7_U377 ( .A(vscale_core_DW01_add_7n102), .ZN(vscale_core_DW01_add_7n100) );
;
  vscale_core_DW01_sub_8 pipeline_md_sub_50_C58 

  XOR2_X2 vscale_core_DW01_sub_8_U1 ( .A(vscale_core_DW01_sub_8n53), .B(vscale_core_DW01_sub_8n1), .Z(pipeline_md_N60) );
  HA_X1 vscale_core_DW01_sub_8_U2 ( .A(vscale_core_DW01_sub_8n54), .B(vscale_core_DW01_sub_8n2), .CO(vscale_core_DW01_sub_8n1), .S(pipeline_md_N59) );
  HA_X1 vscale_core_DW01_sub_8_U3 ( .A(vscale_core_DW01_sub_8n55), .B(vscale_core_DW01_sub_8n3), .CO(vscale_core_DW01_sub_8n2), .S(pipeline_md_N58) );
  HA_X1 vscale_core_DW01_sub_8_U4 ( .A(vscale_core_DW01_sub_8n56), .B(vscale_core_DW01_sub_8n4), .CO(vscale_core_DW01_sub_8n3), .S(pipeline_md_N57) );
  HA_X1 vscale_core_DW01_sub_8_U5 ( .A(vscale_core_DW01_sub_8n57), .B(vscale_core_DW01_sub_8n5), .CO(vscale_core_DW01_sub_8n4), .S(pipeline_md_N56) );
  HA_X1 vscale_core_DW01_sub_8_U6 ( .A(vscale_core_DW01_sub_8n58), .B(vscale_core_DW01_sub_8n6), .CO(vscale_core_DW01_sub_8n5), .S(pipeline_md_N55) );
  HA_X1 vscale_core_DW01_sub_8_U7 ( .A(vscale_core_DW01_sub_8n59), .B(vscale_core_DW01_sub_8n7), .CO(vscale_core_DW01_sub_8n6), .S(pipeline_md_N54) );
  HA_X1 vscale_core_DW01_sub_8_U8 ( .A(vscale_core_DW01_sub_8n60), .B(vscale_core_DW01_sub_8n8), .CO(vscale_core_DW01_sub_8n7), .S(pipeline_md_N53) );
  HA_X1 vscale_core_DW01_sub_8_U9 ( .A(vscale_core_DW01_sub_8n61), .B(vscale_core_DW01_sub_8n9), .CO(vscale_core_DW01_sub_8n8), .S(pipeline_md_N52) );
  HA_X1 vscale_core_DW01_sub_8_U10 ( .A(vscale_core_DW01_sub_8n62), .B(vscale_core_DW01_sub_8n10), .CO(vscale_core_DW01_sub_8n9), .S(pipeline_md_N51) );
  HA_X1 vscale_core_DW01_sub_8_U11 ( .A(vscale_core_DW01_sub_8n63), .B(vscale_core_DW01_sub_8n11), .CO(vscale_core_DW01_sub_8n10), .S(pipeline_md_N50) );
  HA_X1 vscale_core_DW01_sub_8_U12 ( .A(vscale_core_DW01_sub_8n64), .B(vscale_core_DW01_sub_8n12), .CO(vscale_core_DW01_sub_8n11), .S(pipeline_md_N49) );
  HA_X1 vscale_core_DW01_sub_8_U13 ( .A(vscale_core_DW01_sub_8n65), .B(vscale_core_DW01_sub_8n13), .CO(vscale_core_DW01_sub_8n12), .S(pipeline_md_N48) );
  HA_X1 vscale_core_DW01_sub_8_U14 ( .A(vscale_core_DW01_sub_8n66), .B(vscale_core_DW01_sub_8n14), .CO(vscale_core_DW01_sub_8n13), .S(pipeline_md_N47) );
  HA_X1 vscale_core_DW01_sub_8_U15 ( .A(vscale_core_DW01_sub_8n67), .B(vscale_core_DW01_sub_8n15), .CO(vscale_core_DW01_sub_8n14), .S(pipeline_md_N46) );
  HA_X1 vscale_core_DW01_sub_8_U16 ( .A(vscale_core_DW01_sub_8n68), .B(vscale_core_DW01_sub_8n170), .CO(vscale_core_DW01_sub_8n15), .S(pipeline_md_N45) );
  NAND2_X2 vscale_core_DW01_sub_8_U21 ( .A1(vscale_core_DW01_sub_8n24), .A2(vscale_core_DW01_sub_8n19), .ZN(vscale_core_DW01_sub_8n18) );
  XNOR2_X2 vscale_core_DW01_sub_8_U23 ( .A(vscale_core_DW01_sub_8n22), .B(pipeline_rs1_data_bypassed[14]), .ZN(pipeline_md_N43) );
  NAND2_X2 vscale_core_DW01_sub_8_U24 ( .A1(vscale_core_DW01_sub_8n22), .A2(vscale_core_DW01_sub_8n21), .ZN(vscale_core_DW01_sub_8n20) );
  XOR2_X2 vscale_core_DW01_sub_8_U26 ( .A(pipeline_rs1_data_bypassed[13]), .B(vscale_core_DW01_sub_8n25), .Z(pipeline_md_N42) );
  NAND2_X2 vscale_core_DW01_sub_8_U31 ( .A1(vscale_core_DW01_sub_8n28), .A2(vscale_core_DW01_sub_8n26), .ZN(vscale_core_DW01_sub_8n25) );
  NAND2_X2 vscale_core_DW01_sub_8_U36 ( .A1(vscale_core_DW01_sub_8n35), .A2(vscale_core_DW01_sub_8n30), .ZN(vscale_core_DW01_sub_8n29) );
  NAND2_X2 vscale_core_DW01_sub_8_U39 ( .A1(vscale_core_DW01_sub_8n33), .A2(vscale_core_DW01_sub_8n32), .ZN(vscale_core_DW01_sub_8n31) );
  NAND2_X2 vscale_core_DW01_sub_8_U50 ( .A1(vscale_core_DW01_sub_8n43), .A2(vscale_core_DW01_sub_8n40), .ZN(vscale_core_DW01_sub_8n39) );
  NAND2_X2 vscale_core_DW01_sub_8_U55 ( .A1(vscale_core_DW01_sub_8n46), .A2(vscale_core_DW01_sub_8n43), .ZN(vscale_core_DW01_sub_8n42) );
  NAND2_X2 vscale_core_DW01_sub_8_U58 ( .A1(vscale_core_DW01_sub_8n46), .A2(vscale_core_DW01_sub_8n45), .ZN(vscale_core_DW01_sub_8n44) );
  NAND2_X2 vscale_core_DW01_sub_8_U62 ( .A1(vscale_core_DW01_sub_8n48), .A2(vscale_core_DW01_sub_8n51), .ZN(vscale_core_DW01_sub_8n47) );
  BUF_X4 vscale_core_DW01_sub_8_U88 ( .A(pipeline_rs1_data_bypassed[0]), .Z(pipeline_md_N29) );
  XNOR2_X1 vscale_core_DW01_sub_8_U89 ( .A(vscale_core_DW01_sub_8n36), .B(pipeline_rs1_data_bypassed[9]), .ZN(pipeline_md_N38) );
  XOR2_X1 vscale_core_DW01_sub_8_U90 ( .A(pipeline_rs1_data_bypassed[15]), .B(vscale_core_DW01_sub_8n20), .Z(pipeline_md_N44) );
  XNOR2_X1 vscale_core_DW01_sub_8_U91 ( .A(vscale_core_DW01_sub_8n41), .B(pipeline_rs1_data_bypassed[7]), .ZN(pipeline_md_N36) );
  XOR2_X1 vscale_core_DW01_sub_8_U92 ( .A(pipeline_rs1_data_bypassed[0]), .B(n6637), .Z(pipeline_md_N30) );
  INV_X2 vscale_core_DW01_sub_8_U93 ( .A(pipeline_rs1_data_bypassed[27]), .ZN(vscale_core_DW01_sub_8n57) );
  INV_X1 vscale_core_DW01_sub_8_U94 ( .A(pipeline_rs1_data_bypassed[16]), .ZN(vscale_core_DW01_sub_8n68) );
  XNOR2_X1 vscale_core_DW01_sub_8_U95 ( .A(vscale_core_DW01_sub_8n49), .B(pipeline_rs1_data_bypassed[3]), .ZN(pipeline_md_N32) );
  NOR2_X2 vscale_core_DW01_sub_8_U96 ( .A1(vscale_core_DW01_sub_8n37), .A2(vscale_core_DW01_sub_8n29), .ZN(vscale_core_DW01_sub_8n28) );
  NOR2_X2 vscale_core_DW01_sub_8_U97 ( .A1(vscale_core_DW01_sub_8n27), .A2(vscale_core_DW01_sub_8n23), .ZN(vscale_core_DW01_sub_8n22) );
  NOR2_X2 vscale_core_DW01_sub_8_U98 ( .A1(vscale_core_DW01_sub_8n37), .A2(vscale_core_DW01_sub_8n34), .ZN(vscale_core_DW01_sub_8n33) );
  NOR2_X1 vscale_core_DW01_sub_8_U99 ( .A1(n6637), .A2(pipeline_rs1_data_bypassed[0]), .ZN(vscale_core_DW01_sub_8n51) );
  AND2_X1 vscale_core_DW01_sub_8_U100 ( .A1(vscale_core_DW01_sub_8n17), .A2(vscale_core_DW01_sub_8n38), .ZN(vscale_core_DW01_sub_8n170) );
  NOR2_X2 vscale_core_DW01_sub_8_U101 ( .A1(vscale_core_DW01_sub_8n39), .A2(vscale_core_DW01_sub_8n47), .ZN(vscale_core_DW01_sub_8n38) );
  NOR2_X2 vscale_core_DW01_sub_8_U102 ( .A1(vscale_core_DW01_sub_8n29), .A2(vscale_core_DW01_sub_8n18), .ZN(vscale_core_DW01_sub_8n17) );
  NOR2_X1 vscale_core_DW01_sub_8_U103 ( .A1(pipeline_rs1_data_bypassed[14]), .A2(pipeline_rs1_data_bypassed[15]), .ZN(vscale_core_DW01_sub_8n19) );
  NOR2_X1 vscale_core_DW01_sub_8_U104 ( .A1(pipeline_rs1_data_bypassed[12]), .A2(pipeline_rs1_data_bypassed[13]), .ZN(vscale_core_DW01_sub_8n24) );
  XOR2_X1 vscale_core_DW01_sub_8_U105 ( .A(pipeline_rs1_data_bypassed[12]), .B(vscale_core_DW01_sub_8n27), .Z(pipeline_md_N41) );
  INV_X1 vscale_core_DW01_sub_8_U106 ( .A(pipeline_rs1_data_bypassed[12]), .ZN(vscale_core_DW01_sub_8n26) );
  XOR2_X1 vscale_core_DW01_sub_8_U107 ( .A(pipeline_rs1_data_bypassed[11]), .B(vscale_core_DW01_sub_8n31), .Z(pipeline_md_N40) );
  XOR2_X1 vscale_core_DW01_sub_8_U108 ( .A(pipeline_rs1_data_bypassed[5]), .B(vscale_core_DW01_sub_8n44), .Z(pipeline_md_N34) );
  XOR2_X1 vscale_core_DW01_sub_8_U109 ( .A(pipeline_rs1_data_bypassed[6]), .B(vscale_core_DW01_sub_8n42), .Z(pipeline_md_N35) );
  NOR2_X1 vscale_core_DW01_sub_8_U110 ( .A1(vscale_core_DW01_sub_8n42), .A2(pipeline_rs1_data_bypassed[6]), .ZN(vscale_core_DW01_sub_8n41) );
  NOR2_X1 vscale_core_DW01_sub_8_U111 ( .A1(pipeline_rs1_data_bypassed[6]), .A2(pipeline_rs1_data_bypassed[7]), .ZN(vscale_core_DW01_sub_8n40) );
  XOR2_X1 vscale_core_DW01_sub_8_U112 ( .A(pipeline_rs1_data_bypassed[2]), .B(vscale_core_DW01_sub_8n50), .Z(pipeline_md_N31) );
  NOR2_X1 vscale_core_DW01_sub_8_U113 ( .A1(vscale_core_DW01_sub_8n50), .A2(pipeline_rs1_data_bypassed[2]), .ZN(vscale_core_DW01_sub_8n49) );
  NOR2_X1 vscale_core_DW01_sub_8_U114 ( .A1(pipeline_rs1_data_bypassed[2]), .A2(pipeline_rs1_data_bypassed[3]), .ZN(vscale_core_DW01_sub_8n48) );
  XNOR2_X1 vscale_core_DW01_sub_8_U115 ( .A(vscale_core_DW01_sub_8n33), .B(pipeline_rs1_data_bypassed[10]), .ZN(pipeline_md_N39) );
  INV_X2 vscale_core_DW01_sub_8_U116 ( .A(pipeline_rs1_data_bypassed[10]), .ZN(vscale_core_DW01_sub_8n32) );
  NOR2_X1 vscale_core_DW01_sub_8_U117 ( .A1(pipeline_rs1_data_bypassed[10]), .A2(pipeline_rs1_data_bypassed[11]), .ZN(vscale_core_DW01_sub_8n30) );
  XOR2_X1 vscale_core_DW01_sub_8_U118 ( .A(pipeline_rs1_data_bypassed[8]), .B(vscale_core_DW01_sub_8n37), .Z(pipeline_md_N37) );
  NOR2_X1 vscale_core_DW01_sub_8_U119 ( .A1(vscale_core_DW01_sub_8n37), .A2(pipeline_rs1_data_bypassed[8]), .ZN(vscale_core_DW01_sub_8n36) );
  NOR2_X1 vscale_core_DW01_sub_8_U120 ( .A1(pipeline_rs1_data_bypassed[8]), .A2(pipeline_rs1_data_bypassed[9]), .ZN(vscale_core_DW01_sub_8n35) );
  XNOR2_X1 vscale_core_DW01_sub_8_U121 ( .A(vscale_core_DW01_sub_8n46), .B(n6998), .ZN(pipeline_md_N33) );
  INV_X2 vscale_core_DW01_sub_8_U122 ( .A(n6998), .ZN(vscale_core_DW01_sub_8n45) );
  NOR2_X1 vscale_core_DW01_sub_8_U123 ( .A1(n6998), .A2(pipeline_rs1_data_bypassed[5]), .ZN(vscale_core_DW01_sub_8n43) );
  INV_X4 vscale_core_DW01_sub_8_U124 ( .A(pipeline_rs1_data_bypassed[17]), .ZN(vscale_core_DW01_sub_8n67) );
  INV_X4 vscale_core_DW01_sub_8_U125 ( .A(pipeline_rs1_data_bypassed[18]), .ZN(vscale_core_DW01_sub_8n66) );
  INV_X4 vscale_core_DW01_sub_8_U126 ( .A(pipeline_rs1_data_bypassed[19]), .ZN(vscale_core_DW01_sub_8n65) );
  INV_X4 vscale_core_DW01_sub_8_U127 ( .A(pipeline_rs1_data_bypassed[20]), .ZN(vscale_core_DW01_sub_8n64) );
  INV_X4 vscale_core_DW01_sub_8_U128 ( .A(pipeline_rs1_data_bypassed[21]), .ZN(vscale_core_DW01_sub_8n63) );
  INV_X4 vscale_core_DW01_sub_8_U129 ( .A(pipeline_rs1_data_bypassed[22]), .ZN(vscale_core_DW01_sub_8n62) );
  INV_X4 vscale_core_DW01_sub_8_U130 ( .A(n6979), .ZN(vscale_core_DW01_sub_8n61) );
  INV_X4 vscale_core_DW01_sub_8_U131 ( .A(pipeline_rs1_data_bypassed[24]), .ZN(vscale_core_DW01_sub_8n60) );
  INV_X4 vscale_core_DW01_sub_8_U132 ( .A(pipeline_rs1_data_bypassed[25]), .ZN(vscale_core_DW01_sub_8n59) );
  INV_X4 vscale_core_DW01_sub_8_U133 ( .A(pipeline_rs1_data_bypassed[26]), .ZN(vscale_core_DW01_sub_8n58) );
  INV_X4 vscale_core_DW01_sub_8_U134 ( .A(pipeline_rs1_data_bypassed[28]), .ZN(vscale_core_DW01_sub_8n56) );
  INV_X4 vscale_core_DW01_sub_8_U135 ( .A(pipeline_rs1_data_bypassed[29]), .ZN(vscale_core_DW01_sub_8n55) );
  INV_X4 vscale_core_DW01_sub_8_U136 ( .A(pipeline_rs1_data_bypassed[30]), .ZN(vscale_core_DW01_sub_8n54) );
  INV_X4 vscale_core_DW01_sub_8_U137 ( .A(pipeline_rs1_data_bypassed[31]), .ZN(vscale_core_DW01_sub_8n53) );
  INV_X4 vscale_core_DW01_sub_8_U138 ( .A(vscale_core_DW01_sub_8n51), .ZN(vscale_core_DW01_sub_8n50) );
  INV_X4 vscale_core_DW01_sub_8_U139 ( .A(vscale_core_DW01_sub_8n47), .ZN(vscale_core_DW01_sub_8n46) );
  INV_X4 vscale_core_DW01_sub_8_U140 ( .A(vscale_core_DW01_sub_8n38), .ZN(vscale_core_DW01_sub_8n37) );
  INV_X4 vscale_core_DW01_sub_8_U141 ( .A(vscale_core_DW01_sub_8n35), .ZN(vscale_core_DW01_sub_8n34) );
  INV_X4 vscale_core_DW01_sub_8_U142 ( .A(vscale_core_DW01_sub_8n28), .ZN(vscale_core_DW01_sub_8n27) );
  INV_X4 vscale_core_DW01_sub_8_U143 ( .A(vscale_core_DW01_sub_8n24), .ZN(vscale_core_DW01_sub_8n23) );
  INV_X4 vscale_core_DW01_sub_8_U144 ( .A(pipeline_rs1_data_bypassed[14]), .ZN(vscale_core_DW01_sub_8n21) );
;
  vscale_core_DW01_sub_9 pipeline_md_sub_50_C60 

  HA_X1 vscale_core_DW01_sub_9_U2 ( .A(vscale_core_DW01_sub_9n54), .B(vscale_core_DW01_sub_9n2), .CO(vscale_core_DW01_sub_9n1), .S(pipeline_md_N93) );
  HA_X1 vscale_core_DW01_sub_9_U3 ( .A(vscale_core_DW01_sub_9n55), .B(vscale_core_DW01_sub_9n3), .CO(vscale_core_DW01_sub_9n2), .S(pipeline_md_N92) );
  HA_X1 vscale_core_DW01_sub_9_U4 ( .A(vscale_core_DW01_sub_9n56), .B(vscale_core_DW01_sub_9n4), .CO(vscale_core_DW01_sub_9n3), .S(pipeline_md_N91) );
  HA_X1 vscale_core_DW01_sub_9_U5 ( .A(vscale_core_DW01_sub_9n57), .B(vscale_core_DW01_sub_9n5), .CO(vscale_core_DW01_sub_9n4), .S(pipeline_md_N90) );
  HA_X1 vscale_core_DW01_sub_9_U6 ( .A(vscale_core_DW01_sub_9n58), .B(vscale_core_DW01_sub_9n6), .CO(vscale_core_DW01_sub_9n5), .S(pipeline_md_N89) );
  HA_X1 vscale_core_DW01_sub_9_U7 ( .A(vscale_core_DW01_sub_9n59), .B(vscale_core_DW01_sub_9n7), .CO(vscale_core_DW01_sub_9n6), .S(pipeline_md_N88) );
  HA_X1 vscale_core_DW01_sub_9_U8 ( .A(vscale_core_DW01_sub_9n60), .B(vscale_core_DW01_sub_9n8), .CO(vscale_core_DW01_sub_9n7), .S(pipeline_md_N87) );
  HA_X1 vscale_core_DW01_sub_9_U9 ( .A(vscale_core_DW01_sub_9n61), .B(vscale_core_DW01_sub_9n9), .CO(vscale_core_DW01_sub_9n8), .S(pipeline_md_N86) );
  HA_X1 vscale_core_DW01_sub_9_U10 ( .A(vscale_core_DW01_sub_9n62), .B(vscale_core_DW01_sub_9n10), .CO(vscale_core_DW01_sub_9n9), .S(pipeline_md_N85) );
  HA_X1 vscale_core_DW01_sub_9_U11 ( .A(vscale_core_DW01_sub_9n63), .B(vscale_core_DW01_sub_9n11), .CO(vscale_core_DW01_sub_9n10), .S(pipeline_md_N84) );
  HA_X1 vscale_core_DW01_sub_9_U12 ( .A(vscale_core_DW01_sub_9n64), .B(vscale_core_DW01_sub_9n12), .CO(vscale_core_DW01_sub_9n11), .S(pipeline_md_N83) );
  HA_X1 vscale_core_DW01_sub_9_U13 ( .A(vscale_core_DW01_sub_9n65), .B(vscale_core_DW01_sub_9n13), .CO(vscale_core_DW01_sub_9n12), .S(pipeline_md_N82) );
  HA_X1 vscale_core_DW01_sub_9_U14 ( .A(vscale_core_DW01_sub_9n66), .B(vscale_core_DW01_sub_9n14), .CO(vscale_core_DW01_sub_9n13), .S(pipeline_md_N81) );
  HA_X1 vscale_core_DW01_sub_9_U15 ( .A(vscale_core_DW01_sub_9n67), .B(vscale_core_DW01_sub_9n15), .CO(vscale_core_DW01_sub_9n14), .S(pipeline_md_N80) );
  HA_X1 vscale_core_DW01_sub_9_U16 ( .A(vscale_core_DW01_sub_9n68), .B(vscale_core_DW01_sub_9n170), .CO(vscale_core_DW01_sub_9n15), .S(pipeline_md_N79) );
  XOR2_X2 vscale_core_DW01_sub_9_U18 ( .A(pipeline_rs2_data_bypassed[15]), .B(vscale_core_DW01_sub_9n20), .Z(pipeline_md_N78) );
  NAND2_X2 vscale_core_DW01_sub_9_U21 ( .A1(vscale_core_DW01_sub_9n24), .A2(vscale_core_DW01_sub_9n19), .ZN(vscale_core_DW01_sub_9n18) );
  NAND2_X2 vscale_core_DW01_sub_9_U24 ( .A1(vscale_core_DW01_sub_9n22), .A2(vscale_core_DW01_sub_9n21), .ZN(vscale_core_DW01_sub_9n20) );
  XOR2_X2 vscale_core_DW01_sub_9_U26 ( .A(pipeline_rs2_data_bypassed[13]), .B(vscale_core_DW01_sub_9n25), .Z(pipeline_md_N76) );
  NAND2_X2 vscale_core_DW01_sub_9_U31 ( .A1(vscale_core_DW01_sub_9n28), .A2(vscale_core_DW01_sub_9n26), .ZN(vscale_core_DW01_sub_9n25) );
  XOR2_X2 vscale_core_DW01_sub_9_U33 ( .A(pipeline_rs2_data_bypassed[11]), .B(vscale_core_DW01_sub_9n31), .Z(pipeline_md_N74) );
  NAND2_X2 vscale_core_DW01_sub_9_U36 ( .A1(vscale_core_DW01_sub_9n35), .A2(vscale_core_DW01_sub_9n30), .ZN(vscale_core_DW01_sub_9n29) );
  NAND2_X2 vscale_core_DW01_sub_9_U39 ( .A1(vscale_core_DW01_sub_9n33), .A2(vscale_core_DW01_sub_9n32), .ZN(vscale_core_DW01_sub_9n31) );
  XNOR2_X2 vscale_core_DW01_sub_9_U41 ( .A(vscale_core_DW01_sub_9n36), .B(pipeline_rs2_data_bypassed[9]), .ZN(pipeline_md_N72) );
  NAND2_X2 vscale_core_DW01_sub_9_U50 ( .A1(vscale_core_DW01_sub_9n43), .A2(vscale_core_DW01_sub_9n40), .ZN(vscale_core_DW01_sub_9n39) );
  XOR2_X2 vscale_core_DW01_sub_9_U52 ( .A(pipeline_rs2_data_bypassed[6]), .B(vscale_core_DW01_sub_9n42), .Z(pipeline_md_N69) );
  NAND2_X2 vscale_core_DW01_sub_9_U55 ( .A1(vscale_core_DW01_sub_9n46), .A2(vscale_core_DW01_sub_9n43), .ZN(vscale_core_DW01_sub_9n42) );
  NAND2_X2 vscale_core_DW01_sub_9_U58 ( .A1(vscale_core_DW01_sub_9n46), .A2(vscale_core_DW01_sub_9n45), .ZN(vscale_core_DW01_sub_9n44) );
  NAND2_X2 vscale_core_DW01_sub_9_U62 ( .A1(vscale_core_DW01_sub_9n48), .A2(vscale_core_DW01_sub_9n51), .ZN(vscale_core_DW01_sub_9n47) );
  XNOR2_X1 vscale_core_DW01_sub_9_U88 ( .A(vscale_core_DW01_sub_9n22), .B(pipeline_rs2_data_bypassed[14]), .ZN(pipeline_md_N77) );
  INV_X1 vscale_core_DW01_sub_9_U89 ( .A(pipeline_rs2_data_bypassed[14]), .ZN(vscale_core_DW01_sub_9n21) );
  XNOR2_X1 vscale_core_DW01_sub_9_U90 ( .A(vscale_core_DW01_sub_9n33), .B(pipeline_rs2_data_bypassed[10]), .ZN(pipeline_md_N73) );
  INV_X1 vscale_core_DW01_sub_9_U91 ( .A(pipeline_rs2_data_bypassed[10]), .ZN(vscale_core_DW01_sub_9n32) );
  XOR2_X1 vscale_core_DW01_sub_9_U92 ( .A(pipeline_rs2_data_bypassed[2]), .B(vscale_core_DW01_sub_9n50), .Z(pipeline_md_N65) );
  XOR2_X1 vscale_core_DW01_sub_9_U93 ( .A(pipeline_rs2_data_bypassed[5]), .B(vscale_core_DW01_sub_9n44), .Z(pipeline_md_N68) );
  INV_X1 vscale_core_DW01_sub_9_U94 ( .A(pipeline_rs2_data_bypassed[16]), .ZN(vscale_core_DW01_sub_9n68) );
  NOR2_X1 vscale_core_DW01_sub_9_U95 ( .A1(vscale_core_DW01_sub_9n50), .A2(pipeline_rs2_data_bypassed[2]), .ZN(vscale_core_DW01_sub_9n49) );
  XNOR2_X1 vscale_core_DW01_sub_9_U96 ( .A(pipeline_rs2_data_bypassed[31]), .B(vscale_core_DW01_sub_9n1), .ZN(pipeline_md_N94) );
  NOR2_X2 vscale_core_DW01_sub_9_U97 ( .A1(vscale_core_DW01_sub_9n37), .A2(vscale_core_DW01_sub_9n29), .ZN(vscale_core_DW01_sub_9n28) );
  NOR2_X2 vscale_core_DW01_sub_9_U98 ( .A1(vscale_core_DW01_sub_9n37), .A2(vscale_core_DW01_sub_9n34), .ZN(vscale_core_DW01_sub_9n33) );
  NOR2_X2 vscale_core_DW01_sub_9_U99 ( .A1(vscale_core_DW01_sub_9n27), .A2(vscale_core_DW01_sub_9n23), .ZN(vscale_core_DW01_sub_9n22) );
  NOR2_X1 vscale_core_DW01_sub_9_U100 ( .A1(pipeline_rs2_data_bypassed[10]), .A2(pipeline_rs2_data_bypassed[11]), .ZN(vscale_core_DW01_sub_9n30) );
  AND2_X1 vscale_core_DW01_sub_9_U101 ( .A1(vscale_core_DW01_sub_9n17), .A2(vscale_core_DW01_sub_9n38), .ZN(vscale_core_DW01_sub_9n170) );
  NOR2_X2 vscale_core_DW01_sub_9_U102 ( .A1(vscale_core_DW01_sub_9n39), .A2(vscale_core_DW01_sub_9n47), .ZN(vscale_core_DW01_sub_9n38) );
  NOR2_X2 vscale_core_DW01_sub_9_U103 ( .A1(vscale_core_DW01_sub_9n29), .A2(vscale_core_DW01_sub_9n18), .ZN(vscale_core_DW01_sub_9n17) );
  NOR2_X1 vscale_core_DW01_sub_9_U104 ( .A1(pipeline_rs2_data_bypassed[14]), .A2(pipeline_rs2_data_bypassed[15]), .ZN(vscale_core_DW01_sub_9n19) );
  NOR2_X1 vscale_core_DW01_sub_9_U105 ( .A1(vscale_core_DW01_sub_9n42), .A2(pipeline_rs2_data_bypassed[6]), .ZN(vscale_core_DW01_sub_9n41) );
  BUF_X4 vscale_core_DW01_sub_9_U106 ( .A(pipeline_rs2_data_bypassed[0]), .Z(pipeline_md_N63) );
  NOR2_X1 vscale_core_DW01_sub_9_U107 ( .A1(n7004), .A2(pipeline_rs2_data_bypassed[5]), .ZN(vscale_core_DW01_sub_9n43) );
  XNOR2_X1 vscale_core_DW01_sub_9_U108 ( .A(vscale_core_DW01_sub_9n46), .B(n7004), .ZN(pipeline_md_N67) );
  INV_X1 vscale_core_DW01_sub_9_U109 ( .A(n7004), .ZN(vscale_core_DW01_sub_9n45) );
  NOR2_X1 vscale_core_DW01_sub_9_U110 ( .A1(pipeline_rs2_data_bypassed[1]), .A2(pipeline_rs2_data_bypassed[0]), .ZN(vscale_core_DW01_sub_9n51) );
  XOR2_X1 vscale_core_DW01_sub_9_U111 ( .A(pipeline_rs2_data_bypassed[0]), .B(pipeline_rs2_data_bypassed[1]), .Z(pipeline_md_N64) );
  NOR2_X1 vscale_core_DW01_sub_9_U112 ( .A1(pipeline_rs2_data_bypassed[8]), .A2(pipeline_rs2_data_bypassed[9]), .ZN(vscale_core_DW01_sub_9n35) );
  XOR2_X1 vscale_core_DW01_sub_9_U113 ( .A(pipeline_rs2_data_bypassed[8]), .B(vscale_core_DW01_sub_9n37), .Z(pipeline_md_N71) );
  NOR2_X1 vscale_core_DW01_sub_9_U114 ( .A1(vscale_core_DW01_sub_9n37), .A2(pipeline_rs2_data_bypassed[8]), .ZN(vscale_core_DW01_sub_9n36) );
  XOR2_X1 vscale_core_DW01_sub_9_U115 ( .A(pipeline_rs2_data_bypassed[12]), .B(vscale_core_DW01_sub_9n27), .Z(pipeline_md_N75) );
  INV_X2 vscale_core_DW01_sub_9_U116 ( .A(pipeline_rs2_data_bypassed[12]), .ZN(vscale_core_DW01_sub_9n26) );
  NOR2_X1 vscale_core_DW01_sub_9_U117 ( .A1(pipeline_rs2_data_bypassed[12]), .A2(pipeline_rs2_data_bypassed[13]), .ZN(vscale_core_DW01_sub_9n24) );
  XNOR2_X1 vscale_core_DW01_sub_9_U118 ( .A(vscale_core_DW01_sub_9n41), .B(pipeline_rs2_data_bypassed[7]), .ZN(pipeline_md_N70) );
  NOR2_X1 vscale_core_DW01_sub_9_U119 ( .A1(pipeline_rs2_data_bypassed[6]), .A2(pipeline_rs2_data_bypassed[7]), .ZN(vscale_core_DW01_sub_9n40) );
  XNOR2_X1 vscale_core_DW01_sub_9_U120 ( .A(vscale_core_DW01_sub_9n49), .B(n6987), .ZN(pipeline_md_N66) );
  NOR2_X1 vscale_core_DW01_sub_9_U121 ( .A1(pipeline_rs2_data_bypassed[2]), .A2(n6987), .ZN(vscale_core_DW01_sub_9n48) );
  INV_X4 vscale_core_DW01_sub_9_U122 ( .A(pipeline_rs2_data_bypassed[17]), .ZN(vscale_core_DW01_sub_9n67) );
  INV_X4 vscale_core_DW01_sub_9_U123 ( .A(pipeline_rs2_data_bypassed[18]), .ZN(vscale_core_DW01_sub_9n66) );
  INV_X4 vscale_core_DW01_sub_9_U124 ( .A(pipeline_rs2_data_bypassed[19]), .ZN(vscale_core_DW01_sub_9n65) );
  INV_X4 vscale_core_DW01_sub_9_U125 ( .A(pipeline_rs2_data_bypassed[20]), .ZN(vscale_core_DW01_sub_9n64) );
  INV_X4 vscale_core_DW01_sub_9_U126 ( .A(pipeline_rs2_data_bypassed[21]), .ZN(vscale_core_DW01_sub_9n63) );
  INV_X4 vscale_core_DW01_sub_9_U127 ( .A(pipeline_rs2_data_bypassed[22]), .ZN(vscale_core_DW01_sub_9n62) );
  INV_X4 vscale_core_DW01_sub_9_U128 ( .A(pipeline_rs2_data_bypassed[23]), .ZN(vscale_core_DW01_sub_9n61) );
  INV_X4 vscale_core_DW01_sub_9_U129 ( .A(pipeline_rs2_data_bypassed[24]), .ZN(vscale_core_DW01_sub_9n60) );
  INV_X4 vscale_core_DW01_sub_9_U130 ( .A(pipeline_rs2_data_bypassed[25]), .ZN(vscale_core_DW01_sub_9n59) );
  INV_X4 vscale_core_DW01_sub_9_U131 ( .A(pipeline_rs2_data_bypassed[26]), .ZN(vscale_core_DW01_sub_9n58) );
  INV_X4 vscale_core_DW01_sub_9_U132 ( .A(pipeline_rs2_data_bypassed[27]), .ZN(vscale_core_DW01_sub_9n57) );
  INV_X4 vscale_core_DW01_sub_9_U133 ( .A(pipeline_rs2_data_bypassed[28]), .ZN(vscale_core_DW01_sub_9n56) );
  INV_X4 vscale_core_DW01_sub_9_U134 ( .A(pipeline_rs2_data_bypassed[29]), .ZN(vscale_core_DW01_sub_9n55) );
  INV_X4 vscale_core_DW01_sub_9_U135 ( .A(pipeline_rs2_data_bypassed[30]), .ZN(vscale_core_DW01_sub_9n54) );
  INV_X4 vscale_core_DW01_sub_9_U136 ( .A(vscale_core_DW01_sub_9n51), .ZN(vscale_core_DW01_sub_9n50) );
  INV_X4 vscale_core_DW01_sub_9_U137 ( .A(vscale_core_DW01_sub_9n47), .ZN(vscale_core_DW01_sub_9n46) );
  INV_X4 vscale_core_DW01_sub_9_U138 ( .A(vscale_core_DW01_sub_9n38), .ZN(vscale_core_DW01_sub_9n37) );
  INV_X4 vscale_core_DW01_sub_9_U139 ( .A(vscale_core_DW01_sub_9n35), .ZN(vscale_core_DW01_sub_9n34) );
  INV_X4 vscale_core_DW01_sub_9_U140 ( .A(vscale_core_DW01_sub_9n28), .ZN(vscale_core_DW01_sub_9n27) );
  INV_X4 vscale_core_DW01_sub_9_U141 ( .A(vscale_core_DW01_sub_9n24), .ZN(vscale_core_DW01_sub_9n23) );
;
  vscale_core_DW01_inc_4 pipeline_csr_add_314 

  XOR2_X2 vscale_core_DW01_inc_4_U1 ( .A(pipeline_csr_instret_full[63]), .B(vscale_core_DW01_inc_4n1), .Z(pipeline_csr_N839) );
  HA_X1 vscale_core_DW01_inc_4_U2 ( .A(pipeline_csr_instret_full[62]), .B(vscale_core_DW01_inc_4n2), .CO(vscale_core_DW01_inc_4n1), .S(pipeline_csr_N838) );
  HA_X1 vscale_core_DW01_inc_4_U3 ( .A(pipeline_csr_instret_full[61]), .B(vscale_core_DW01_inc_4n3), .CO(vscale_core_DW01_inc_4n2), .S(pipeline_csr_N837) );
  HA_X1 vscale_core_DW01_inc_4_U4 ( .A(pipeline_csr_instret_full[60]), .B(vscale_core_DW01_inc_4n4), .CO(vscale_core_DW01_inc_4n3), .S(pipeline_csr_N836) );
  HA_X1 vscale_core_DW01_inc_4_U5 ( .A(pipeline_csr_instret_full[59]), .B(vscale_core_DW01_inc_4n5), .CO(vscale_core_DW01_inc_4n4), .S(pipeline_csr_N835) );
  HA_X1 vscale_core_DW01_inc_4_U6 ( .A(pipeline_csr_instret_full[58]), .B(vscale_core_DW01_inc_4n6), .CO(vscale_core_DW01_inc_4n5), .S(pipeline_csr_N834) );
  HA_X1 vscale_core_DW01_inc_4_U7 ( .A(pipeline_csr_instret_full[57]), .B(vscale_core_DW01_inc_4n7), .CO(vscale_core_DW01_inc_4n6), .S(pipeline_csr_N833) );
  HA_X1 vscale_core_DW01_inc_4_U8 ( .A(pipeline_csr_instret_full[56]), .B(vscale_core_DW01_inc_4n8), .CO(vscale_core_DW01_inc_4n7), .S(pipeline_csr_N832) );
  HA_X1 vscale_core_DW01_inc_4_U9 ( .A(pipeline_csr_instret_full[55]), .B(vscale_core_DW01_inc_4n9), .CO(vscale_core_DW01_inc_4n8), .S(pipeline_csr_N831) );
  HA_X1 vscale_core_DW01_inc_4_U10 ( .A(pipeline_csr_instret_full[54]), .B(vscale_core_DW01_inc_4n10), .CO(vscale_core_DW01_inc_4n9), .S(pipeline_csr_N830) );
  HA_X1 vscale_core_DW01_inc_4_U11 ( .A(pipeline_csr_instret_full[53]), .B(vscale_core_DW01_inc_4n11), .CO(vscale_core_DW01_inc_4n10), .S(pipeline_csr_N829) );
  HA_X1 vscale_core_DW01_inc_4_U12 ( .A(n10889), .B(vscale_core_DW01_inc_4n12), .CO(vscale_core_DW01_inc_4n11), .S(pipeline_csr_N828) );
  HA_X1 vscale_core_DW01_inc_4_U13 ( .A(pipeline_csr_instret_full[51]), .B(vscale_core_DW01_inc_4n13), .CO(vscale_core_DW01_inc_4n12), .S(pipeline_csr_N827) );
  HA_X1 vscale_core_DW01_inc_4_U14 ( .A(pipeline_csr_instret_full[50]), .B(vscale_core_DW01_inc_4n14), .CO(vscale_core_DW01_inc_4n13), .S(pipeline_csr_N826) );
  HA_X1 vscale_core_DW01_inc_4_U15 ( .A(pipeline_csr_instret_full[49]), .B(vscale_core_DW01_inc_4n15), .CO(vscale_core_DW01_inc_4n14), .S(pipeline_csr_N825) );
  HA_X1 vscale_core_DW01_inc_4_U16 ( .A(pipeline_csr_instret_full[48]), .B(vscale_core_DW01_inc_4n16), .CO(vscale_core_DW01_inc_4n15), .S(pipeline_csr_N824) );
  HA_X1 vscale_core_DW01_inc_4_U17 ( .A(n11104), .B(vscale_core_DW01_inc_4n17), .CO(vscale_core_DW01_inc_4n16), .S(pipeline_csr_N823) );
  HA_X1 vscale_core_DW01_inc_4_U18 ( .A(pipeline_csr_instret_full[46]), .B(vscale_core_DW01_inc_4n18), .CO(vscale_core_DW01_inc_4n17), .S(pipeline_csr_N822) );
  HA_X1 vscale_core_DW01_inc_4_U19 ( .A(pipeline_csr_instret_full[45]), .B(vscale_core_DW01_inc_4n19), .CO(vscale_core_DW01_inc_4n18), .S(pipeline_csr_N821) );
  HA_X1 vscale_core_DW01_inc_4_U20 ( .A(pipeline_csr_instret_full[44]), .B(vscale_core_DW01_inc_4n20), .CO(vscale_core_DW01_inc_4n19), .S(pipeline_csr_N820) );
  HA_X1 vscale_core_DW01_inc_4_U21 ( .A(pipeline_csr_instret_full[43]), .B(vscale_core_DW01_inc_4n21), .CO(vscale_core_DW01_inc_4n20), .S(pipeline_csr_N819) );
  HA_X1 vscale_core_DW01_inc_4_U22 ( .A(pipeline_csr_instret_full[42]), .B(vscale_core_DW01_inc_4n22), .CO(vscale_core_DW01_inc_4n21), .S(pipeline_csr_N818) );
  XOR2_X2 vscale_core_DW01_inc_4_U23 ( .A(vscale_core_DW01_inc_4n25), .B(vscale_core_DW01_inc_4n26), .Z(pipeline_csr_N817) );
  NAND2_X2 vscale_core_DW01_inc_4_U25 ( .A1(vscale_core_DW01_inc_4n27), .A2(pipeline_csr_instret_full[41]), .ZN(vscale_core_DW01_inc_4n23) );
  XOR2_X2 vscale_core_DW01_inc_4_U28 ( .A(vscale_core_DW01_inc_4n28), .B(vscale_core_DW01_inc_4n29), .Z(pipeline_csr_N816) );
  NAND2_X2 vscale_core_DW01_inc_4_U29 ( .A1(vscale_core_DW01_inc_4n67), .A2(vscale_core_DW01_inc_4n27), .ZN(vscale_core_DW01_inc_4n26) );
  XNOR2_X2 vscale_core_DW01_inc_4_U32 ( .A(vscale_core_DW01_inc_4n36), .B(vscale_core_DW01_inc_4n35), .ZN(pipeline_csr_N815) );
  NAND2_X2 vscale_core_DW01_inc_4_U33 ( .A1(vscale_core_DW01_inc_4n67), .A2(vscale_core_DW01_inc_4n30), .ZN(vscale_core_DW01_inc_4n29) );
  NAND2_X2 vscale_core_DW01_inc_4_U35 ( .A1(vscale_core_DW01_inc_4n51), .A2(vscale_core_DW01_inc_4n32), .ZN(vscale_core_DW01_inc_4n31) );
  NAND2_X2 vscale_core_DW01_inc_4_U37 ( .A1(pipeline_csr_instret_full[38]), .A2(pipeline_csr_instret_full[39]), .ZN(vscale_core_DW01_inc_4n33) );
  XOR2_X2 vscale_core_DW01_inc_4_U40 ( .A(vscale_core_DW01_inc_4n39), .B(vscale_core_DW01_inc_4n40), .Z(pipeline_csr_N814) );
  XNOR2_X2 vscale_core_DW01_inc_4_U45 ( .A(vscale_core_DW01_inc_4n45), .B(vscale_core_DW01_inc_4n44), .ZN(pipeline_csr_N813) );
  NAND2_X2 vscale_core_DW01_inc_4_U46 ( .A1(vscale_core_DW01_inc_4n49), .A2(vscale_core_DW01_inc_4n41), .ZN(vscale_core_DW01_inc_4n40) );
  NAND2_X2 vscale_core_DW01_inc_4_U48 ( .A1(pipeline_csr_instret_full[36]), .A2(pipeline_csr_instret_full[37]), .ZN(vscale_core_DW01_inc_4n42) );
  XNOR2_X2 vscale_core_DW01_inc_4_U51 ( .A(vscale_core_DW01_inc_4n49), .B(vscale_core_DW01_inc_4n48), .ZN(pipeline_csr_N812) );
  XNOR2_X2 vscale_core_DW01_inc_4_U56 ( .A(vscale_core_DW01_inc_4n55), .B(vscale_core_DW01_inc_4n54), .ZN(pipeline_csr_N811) );
  NAND2_X2 vscale_core_DW01_inc_4_U58 ( .A1(vscale_core_DW01_inc_4n67), .A2(vscale_core_DW01_inc_4n51), .ZN(vscale_core_DW01_inc_4n50) );
  NAND2_X2 vscale_core_DW01_inc_4_U60 ( .A1(pipeline_csr_instret_full[34]), .A2(pipeline_csr_instret_full[35]), .ZN(vscale_core_DW01_inc_4n52) );
  XOR2_X2 vscale_core_DW01_inc_4_U63 ( .A(vscale_core_DW01_inc_4n58), .B(vscale_core_DW01_inc_4n59), .Z(pipeline_csr_N810) );
  XOR2_X2 vscale_core_DW01_inc_4_U68 ( .A(vscale_core_DW01_inc_4n63), .B(vscale_core_DW01_inc_4n64), .Z(pipeline_csr_N809) );
  NAND2_X2 vscale_core_DW01_inc_4_U69 ( .A1(vscale_core_DW01_inc_4n67), .A2(vscale_core_DW01_inc_4n60), .ZN(vscale_core_DW01_inc_4n59) );
  NAND2_X2 vscale_core_DW01_inc_4_U71 ( .A1(pipeline_csr_instret_full[32]), .A2(pipeline_csr_instret_full[33]), .ZN(vscale_core_DW01_inc_4n61) );
  XNOR2_X2 vscale_core_DW01_inc_4_U74 ( .A(vscale_core_DW01_inc_4n67), .B(vscale_core_DW01_inc_4n66), .ZN(pipeline_csr_N808) );
  NAND2_X2 vscale_core_DW01_inc_4_U75 ( .A1(vscale_core_DW01_inc_4n67), .A2(pipeline_csr_instret_full[32]), .ZN(vscale_core_DW01_inc_4n64) );
  XOR2_X2 vscale_core_DW01_inc_4_U78 ( .A(vscale_core_DW01_inc_4n74), .B(vscale_core_DW01_inc_4n75), .Z(pipeline_csr_N807) );
  NAND2_X2 vscale_core_DW01_inc_4_U80 ( .A1(vscale_core_DW01_inc_4n69), .A2(vscale_core_DW01_inc_4n138), .ZN(vscale_core_DW01_inc_4n68) );
  NAND2_X2 vscale_core_DW01_inc_4_U82 ( .A1(vscale_core_DW01_inc_4n88), .A2(vscale_core_DW01_inc_4n71), .ZN(vscale_core_DW01_inc_4n70) );
  NAND2_X2 vscale_core_DW01_inc_4_U84 ( .A1(pipeline_csr_instret_full[30]), .A2(pipeline_csr_instret_full[31]), .ZN(vscale_core_DW01_inc_4n72) );
  XNOR2_X2 vscale_core_DW01_inc_4_U87 ( .A(vscale_core_DW01_inc_4n78), .B(vscale_core_DW01_inc_4n77), .ZN(pipeline_csr_N806) );
  NAND2_X2 vscale_core_DW01_inc_4_U88 ( .A1(vscale_core_DW01_inc_4n78), .A2(pipeline_csr_instret_full[30]), .ZN(vscale_core_DW01_inc_4n75) );
  XOR2_X2 vscale_core_DW01_inc_4_U91 ( .A(vscale_core_DW01_inc_4n81), .B(vscale_core_DW01_inc_4n82), .Z(pipeline_csr_N805) );
  NAND2_X2 vscale_core_DW01_inc_4_U93 ( .A1(pipeline_csr_instret_full[28]), .A2(pipeline_csr_instret_full[29]), .ZN(vscale_core_DW01_inc_4n79) );
  XOR2_X2 vscale_core_DW01_inc_4_U96 ( .A(vscale_core_DW01_inc_4n84), .B(vscale_core_DW01_inc_4n85), .Z(pipeline_csr_N804) );
  NAND2_X2 vscale_core_DW01_inc_4_U97 ( .A1(vscale_core_DW01_inc_4n86), .A2(pipeline_csr_instret_full[28]), .ZN(vscale_core_DW01_inc_4n82) );
  XOR2_X2 vscale_core_DW01_inc_4_U100 ( .A(vscale_core_DW01_inc_4n91), .B(vscale_core_DW01_inc_4n92), .Z(pipeline_csr_N803) );
  NAND2_X2 vscale_core_DW01_inc_4_U105 ( .A1(pipeline_csr_instret_full[26]), .A2(pipeline_csr_instret_full[27]), .ZN(vscale_core_DW01_inc_4n89) );
  XNOR2_X2 vscale_core_DW01_inc_4_U108 ( .A(vscale_core_DW01_inc_4n95), .B(vscale_core_DW01_inc_4n94), .ZN(pipeline_csr_N802) );
  NAND2_X2 vscale_core_DW01_inc_4_U109 ( .A1(vscale_core_DW01_inc_4n95), .A2(pipeline_csr_instret_full[26]), .ZN(vscale_core_DW01_inc_4n92) );
  XOR2_X2 vscale_core_DW01_inc_4_U112 ( .A(vscale_core_DW01_inc_4n98), .B(vscale_core_DW01_inc_4n99), .Z(pipeline_csr_N801) );
  NAND2_X2 vscale_core_DW01_inc_4_U114 ( .A1(pipeline_csr_instret_full[24]), .A2(pipeline_csr_instret_full[25]), .ZN(vscale_core_DW01_inc_4n96) );
  XOR2_X2 vscale_core_DW01_inc_4_U117 ( .A(vscale_core_DW01_inc_4n101), .B(vscale_core_DW01_inc_4n102), .Z(pipeline_csr_N800) );
  NAND2_X2 vscale_core_DW01_inc_4_U118 ( .A1(vscale_core_DW01_inc_4n103), .A2(pipeline_csr_instret_full[24]), .ZN(vscale_core_DW01_inc_4n99) );
  XOR2_X2 vscale_core_DW01_inc_4_U121 ( .A(vscale_core_DW01_inc_4n108), .B(vscale_core_DW01_inc_4n109), .Z(pipeline_csr_N799) );
  NAND2_X2 vscale_core_DW01_inc_4_U124 ( .A1(vscale_core_DW01_inc_4n122), .A2(vscale_core_DW01_inc_4n105), .ZN(vscale_core_DW01_inc_4n104) );
  NAND2_X2 vscale_core_DW01_inc_4_U126 ( .A1(pipeline_csr_instret_full[22]), .A2(pipeline_csr_instret_full[23]), .ZN(vscale_core_DW01_inc_4n106) );
  XNOR2_X2 vscale_core_DW01_inc_4_U129 ( .A(vscale_core_DW01_inc_4n112), .B(vscale_core_DW01_inc_4n111), .ZN(pipeline_csr_N798) );
  NAND2_X2 vscale_core_DW01_inc_4_U130 ( .A1(vscale_core_DW01_inc_4n112), .A2(pipeline_csr_instret_full[22]), .ZN(vscale_core_DW01_inc_4n109) );
  XOR2_X2 vscale_core_DW01_inc_4_U133 ( .A(vscale_core_DW01_inc_4n115), .B(vscale_core_DW01_inc_4n116), .Z(pipeline_csr_N797) );
  NAND2_X2 vscale_core_DW01_inc_4_U135 ( .A1(pipeline_csr_instret_full[20]), .A2(pipeline_csr_instret_full[21]), .ZN(vscale_core_DW01_inc_4n113) );
  XOR2_X2 vscale_core_DW01_inc_4_U138 ( .A(vscale_core_DW01_inc_4n118), .B(vscale_core_DW01_inc_4n119), .Z(pipeline_csr_N796) );
  NAND2_X2 vscale_core_DW01_inc_4_U139 ( .A1(vscale_core_DW01_inc_4n120), .A2(pipeline_csr_instret_full[20]), .ZN(vscale_core_DW01_inc_4n116) );
  XOR2_X2 vscale_core_DW01_inc_4_U142 ( .A(vscale_core_DW01_inc_4n125), .B(vscale_core_DW01_inc_4n126), .Z(pipeline_csr_N795) );
  NAND2_X2 vscale_core_DW01_inc_4_U147 ( .A1(pipeline_csr_instret_full[18]), .A2(pipeline_csr_instret_full[19]), .ZN(vscale_core_DW01_inc_4n123) );
  XNOR2_X2 vscale_core_DW01_inc_4_U150 ( .A(vscale_core_DW01_inc_4n129), .B(vscale_core_DW01_inc_4n128), .ZN(pipeline_csr_N794) );
  NAND2_X2 vscale_core_DW01_inc_4_U151 ( .A1(vscale_core_DW01_inc_4n129), .A2(pipeline_csr_instret_full[18]), .ZN(vscale_core_DW01_inc_4n126) );
  XNOR2_X2 vscale_core_DW01_inc_4_U154 ( .A(vscale_core_DW01_inc_4n133), .B(vscale_core_DW01_inc_4n132), .ZN(pipeline_csr_N793) );
  NAND2_X2 vscale_core_DW01_inc_4_U156 ( .A1(pipeline_csr_instret_full[16]), .A2(pipeline_csr_instret_full[17]), .ZN(vscale_core_DW01_inc_4n130) );
  XOR2_X2 vscale_core_DW01_inc_4_U159 ( .A(vscale_core_DW01_inc_4n136), .B(vscale_core_DW01_inc_4n137), .Z(pipeline_csr_N792) );
  XNOR2_X2 vscale_core_DW01_inc_4_U164 ( .A(vscale_core_DW01_inc_4n144), .B(vscale_core_DW01_inc_4n143), .ZN(pipeline_csr_N791) );
  NAND2_X2 vscale_core_DW01_inc_4_U167 ( .A1(vscale_core_DW01_inc_4n159), .A2(vscale_core_DW01_inc_4n140), .ZN(vscale_core_DW01_inc_4n139) );
  NAND2_X2 vscale_core_DW01_inc_4_U169 ( .A1(pipeline_csr_instret_full[14]), .A2(pipeline_csr_instret_full[15]), .ZN(vscale_core_DW01_inc_4n141) );
  XOR2_X2 vscale_core_DW01_inc_4_U172 ( .A(vscale_core_DW01_inc_4n147), .B(vscale_core_DW01_inc_4n148), .Z(pipeline_csr_N790) );
  XNOR2_X2 vscale_core_DW01_inc_4_U177 ( .A(vscale_core_DW01_inc_4n153), .B(vscale_core_DW01_inc_4n152), .ZN(pipeline_csr_N789) );
  NAND2_X2 vscale_core_DW01_inc_4_U178 ( .A1(vscale_core_DW01_inc_4n157), .A2(vscale_core_DW01_inc_4n149), .ZN(vscale_core_DW01_inc_4n148) );
  NAND2_X2 vscale_core_DW01_inc_4_U180 ( .A1(pipeline_csr_instret_full[12]), .A2(pipeline_csr_instret_full[13]), .ZN(vscale_core_DW01_inc_4n150) );
  XNOR2_X2 vscale_core_DW01_inc_4_U183 ( .A(vscale_core_DW01_inc_4n157), .B(vscale_core_DW01_inc_4n156), .ZN(pipeline_csr_N788) );
  XNOR2_X2 vscale_core_DW01_inc_4_U188 ( .A(vscale_core_DW01_inc_4n163), .B(vscale_core_DW01_inc_4n162), .ZN(pipeline_csr_N787) );
  NAND2_X2 vscale_core_DW01_inc_4_U190 ( .A1(vscale_core_DW01_inc_4n175), .A2(vscale_core_DW01_inc_4n159), .ZN(vscale_core_DW01_inc_4n158) );
  NAND2_X2 vscale_core_DW01_inc_4_U192 ( .A1(pipeline_csr_instret_full[10]), .A2(pipeline_csr_instret_full[11]), .ZN(vscale_core_DW01_inc_4n160) );
  XOR2_X2 vscale_core_DW01_inc_4_U195 ( .A(vscale_core_DW01_inc_4n166), .B(vscale_core_DW01_inc_4n167), .Z(pipeline_csr_N786) );
  XOR2_X2 vscale_core_DW01_inc_4_U200 ( .A(vscale_core_DW01_inc_4n171), .B(vscale_core_DW01_inc_4n172), .Z(pipeline_csr_N785) );
  NAND2_X2 vscale_core_DW01_inc_4_U201 ( .A1(vscale_core_DW01_inc_4n175), .A2(vscale_core_DW01_inc_4n168), .ZN(vscale_core_DW01_inc_4n167) );
  NAND2_X2 vscale_core_DW01_inc_4_U203 ( .A1(pipeline_csr_instret_full[8]), .A2(pipeline_csr_instret_full[9]), .ZN(vscale_core_DW01_inc_4n169) );
  XNOR2_X2 vscale_core_DW01_inc_4_U206 ( .A(vscale_core_DW01_inc_4n175), .B(vscale_core_DW01_inc_4n174), .ZN(pipeline_csr_N784) );
  NAND2_X2 vscale_core_DW01_inc_4_U207 ( .A1(vscale_core_DW01_inc_4n175), .A2(pipeline_csr_instret_full[8]), .ZN(vscale_core_DW01_inc_4n172) );
  XOR2_X2 vscale_core_DW01_inc_4_U210 ( .A(vscale_core_DW01_inc_4n180), .B(vscale_core_DW01_inc_4n181), .Z(pipeline_csr_N783) );
  NAND2_X2 vscale_core_DW01_inc_4_U212 ( .A1(vscale_core_DW01_inc_4n177), .A2(vscale_core_DW01_inc_4n193), .ZN(vscale_core_DW01_inc_4n176) );
  NAND2_X2 vscale_core_DW01_inc_4_U214 ( .A1(pipeline_csr_instret_full[6]), .A2(pipeline_csr_instret_full[7]), .ZN(vscale_core_DW01_inc_4n178) );
  XNOR2_X2 vscale_core_DW01_inc_4_U217 ( .A(vscale_core_DW01_inc_4n184), .B(vscale_core_DW01_inc_4n183), .ZN(pipeline_csr_N782) );
  NAND2_X2 vscale_core_DW01_inc_4_U218 ( .A1(vscale_core_DW01_inc_4n184), .A2(pipeline_csr_instret_full[6]), .ZN(vscale_core_DW01_inc_4n181) );
  XNOR2_X2 vscale_core_DW01_inc_4_U221 ( .A(vscale_core_DW01_inc_4n188), .B(vscale_core_DW01_inc_4n187), .ZN(pipeline_csr_N781) );
  NAND2_X2 vscale_core_DW01_inc_4_U223 ( .A1(pipeline_csr_instret_full[4]), .A2(pipeline_csr_instret_full[5]), .ZN(vscale_core_DW01_inc_4n185) );
  XOR2_X2 vscale_core_DW01_inc_4_U226 ( .A(vscale_core_DW01_inc_4n191), .B(vscale_core_DW01_inc_4n192), .Z(pipeline_csr_N780) );
  XOR2_X2 vscale_core_DW01_inc_4_U231 ( .A(vscale_core_DW01_inc_4n196), .B(vscale_core_DW01_inc_4n197), .Z(pipeline_csr_N779) );
  NAND2_X2 vscale_core_DW01_inc_4_U234 ( .A1(pipeline_csr_instret_full[2]), .A2(pipeline_csr_instret_full[3]), .ZN(vscale_core_DW01_inc_4n194) );
  XNOR2_X2 vscale_core_DW01_inc_4_U237 ( .A(vscale_core_DW01_inc_4n200), .B(vscale_core_DW01_inc_4n199), .ZN(pipeline_csr_N778) );
  NAND2_X2 vscale_core_DW01_inc_4_U238 ( .A1(vscale_core_DW01_inc_4n200), .A2(pipeline_csr_instret_full[2]), .ZN(vscale_core_DW01_inc_4n197) );
  XNOR2_X2 vscale_core_DW01_inc_4_U241 ( .A(vscale_core_DW01_inc_4n203), .B(pipeline_csr_instret_full[0]), .ZN(pipeline_csr_N777) );
  NAND2_X2 vscale_core_DW01_inc_4_U243 ( .A1(pipeline_csr_instret_full[1]), .A2(pipeline_csr_instret_full[0]), .ZN(vscale_core_DW01_inc_4n201) );
  NOR2_X2 vscale_core_DW01_inc_4_U248 ( .A1(vscale_core_DW01_inc_4n104), .A2(vscale_core_DW01_inc_4n70), .ZN(vscale_core_DW01_inc_4n69) );
  NOR2_X2 vscale_core_DW01_inc_4_U249 ( .A1(vscale_core_DW01_inc_4n79), .A2(vscale_core_DW01_inc_4n72), .ZN(vscale_core_DW01_inc_4n71) );
  NOR2_X2 vscale_core_DW01_inc_4_U250 ( .A1(vscale_core_DW01_inc_4n31), .A2(vscale_core_DW01_inc_4n28), .ZN(vscale_core_DW01_inc_4n27) );
  NOR2_X2 vscale_core_DW01_inc_4_U251 ( .A1(vscale_core_DW01_inc_4n137), .A2(vscale_core_DW01_inc_4n104), .ZN(vscale_core_DW01_inc_4n103) );
  NOR2_X2 vscale_core_DW01_inc_4_U252 ( .A1(vscale_core_DW01_inc_4n137), .A2(vscale_core_DW01_inc_4n121), .ZN(vscale_core_DW01_inc_4n120) );
  NOR2_X2 vscale_core_DW01_inc_4_U253 ( .A1(vscale_core_DW01_inc_4n102), .A2(vscale_core_DW01_inc_4n87), .ZN(vscale_core_DW01_inc_4n86) );
  NOR2_X2 vscale_core_DW01_inc_4_U254 ( .A1(vscale_core_DW01_inc_4n85), .A2(vscale_core_DW01_inc_4n79), .ZN(vscale_core_DW01_inc_4n78) );
  NOR2_X2 vscale_core_DW01_inc_4_U255 ( .A1(vscale_core_DW01_inc_4n102), .A2(vscale_core_DW01_inc_4n96), .ZN(vscale_core_DW01_inc_4n95) );
  NOR2_X2 vscale_core_DW01_inc_4_U256 ( .A1(vscale_core_DW01_inc_4n119), .A2(vscale_core_DW01_inc_4n113), .ZN(vscale_core_DW01_inc_4n112) );
  NOR2_X2 vscale_core_DW01_inc_4_U257 ( .A1(vscale_core_DW01_inc_4n137), .A2(vscale_core_DW01_inc_4n130), .ZN(vscale_core_DW01_inc_4n129) );
  NOR2_X2 vscale_core_DW01_inc_4_U258 ( .A1(vscale_core_DW01_inc_4n192), .A2(vscale_core_DW01_inc_4n185), .ZN(vscale_core_DW01_inc_4n184) );
  NOR2_X2 vscale_core_DW01_inc_4_U259 ( .A1(vscale_core_DW01_inc_4n137), .A2(vscale_core_DW01_inc_4n136), .ZN(vscale_core_DW01_inc_4n133) );
  NOR2_X2 vscale_core_DW01_inc_4_U260 ( .A1(vscale_core_DW01_inc_4n148), .A2(vscale_core_DW01_inc_4n147), .ZN(vscale_core_DW01_inc_4n144) );
  NOR2_X2 vscale_core_DW01_inc_4_U261 ( .A1(vscale_core_DW01_inc_4n158), .A2(vscale_core_DW01_inc_4n156), .ZN(vscale_core_DW01_inc_4n153) );
  NOR2_X2 vscale_core_DW01_inc_4_U262 ( .A1(vscale_core_DW01_inc_4n167), .A2(vscale_core_DW01_inc_4n166), .ZN(vscale_core_DW01_inc_4n163) );
  NOR2_X2 vscale_core_DW01_inc_4_U263 ( .A1(vscale_core_DW01_inc_4n50), .A2(vscale_core_DW01_inc_4n48), .ZN(vscale_core_DW01_inc_4n45) );
  NOR2_X2 vscale_core_DW01_inc_4_U264 ( .A1(vscale_core_DW01_inc_4n40), .A2(vscale_core_DW01_inc_4n39), .ZN(vscale_core_DW01_inc_4n36) );
  NOR2_X2 vscale_core_DW01_inc_4_U265 ( .A1(vscale_core_DW01_inc_4n59), .A2(vscale_core_DW01_inc_4n58), .ZN(vscale_core_DW01_inc_4n55) );
  NOR2_X2 vscale_core_DW01_inc_4_U266 ( .A1(vscale_core_DW01_inc_4n192), .A2(vscale_core_DW01_inc_4n191), .ZN(vscale_core_DW01_inc_4n188) );
  NOR2_X2 vscale_core_DW01_inc_4_U267 ( .A1(vscale_core_DW01_inc_4n113), .A2(vscale_core_DW01_inc_4n106), .ZN(vscale_core_DW01_inc_4n105) );
  NOR2_X2 vscale_core_DW01_inc_4_U268 ( .A1(vscale_core_DW01_inc_4n42), .A2(vscale_core_DW01_inc_4n33), .ZN(vscale_core_DW01_inc_4n32) );
  NOR2_X2 vscale_core_DW01_inc_4_U269 ( .A1(vscale_core_DW01_inc_4n185), .A2(vscale_core_DW01_inc_4n178), .ZN(vscale_core_DW01_inc_4n177) );
  NOR2_X2 vscale_core_DW01_inc_4_U270 ( .A1(vscale_core_DW01_inc_4n68), .A2(vscale_core_DW01_inc_4n23), .ZN(vscale_core_DW01_inc_4n22) );
  NOR2_X2 vscale_core_DW01_inc_4_U271 ( .A1(vscale_core_DW01_inc_4n130), .A2(vscale_core_DW01_inc_4n123), .ZN(vscale_core_DW01_inc_4n122) );
  NOR2_X2 vscale_core_DW01_inc_4_U272 ( .A1(vscale_core_DW01_inc_4n96), .A2(vscale_core_DW01_inc_4n89), .ZN(vscale_core_DW01_inc_4n88) );
  NOR2_X2 vscale_core_DW01_inc_4_U273 ( .A1(vscale_core_DW01_inc_4n194), .A2(vscale_core_DW01_inc_4n201), .ZN(vscale_core_DW01_inc_4n193) );
  NOR2_X2 vscale_core_DW01_inc_4_U274 ( .A1(vscale_core_DW01_inc_4n139), .A2(vscale_core_DW01_inc_4n176), .ZN(vscale_core_DW01_inc_4n138) );
  NOR2_X2 vscale_core_DW01_inc_4_U275 ( .A1(vscale_core_DW01_inc_4n150), .A2(vscale_core_DW01_inc_4n141), .ZN(vscale_core_DW01_inc_4n140) );
  NOR2_X2 vscale_core_DW01_inc_4_U276 ( .A1(vscale_core_DW01_inc_4n169), .A2(vscale_core_DW01_inc_4n160), .ZN(vscale_core_DW01_inc_4n159) );
  NOR2_X2 vscale_core_DW01_inc_4_U277 ( .A1(vscale_core_DW01_inc_4n61), .A2(vscale_core_DW01_inc_4n52), .ZN(vscale_core_DW01_inc_4n51) );
  INV_X4 vscale_core_DW01_inc_4_U278 ( .A(pipeline_csr_instret_full[25]), .ZN(vscale_core_DW01_inc_4n98) );
  INV_X4 vscale_core_DW01_inc_4_U279 ( .A(pipeline_csr_instret_full[26]), .ZN(vscale_core_DW01_inc_4n94) );
  INV_X4 vscale_core_DW01_inc_4_U280 ( .A(pipeline_csr_instret_full[27]), .ZN(vscale_core_DW01_inc_4n91) );
  INV_X4 vscale_core_DW01_inc_4_U281 ( .A(vscale_core_DW01_inc_4n88), .ZN(vscale_core_DW01_inc_4n87) );
  INV_X4 vscale_core_DW01_inc_4_U282 ( .A(vscale_core_DW01_inc_4n86), .ZN(vscale_core_DW01_inc_4n85) );
  INV_X4 vscale_core_DW01_inc_4_U283 ( .A(pipeline_csr_instret_full[28]), .ZN(vscale_core_DW01_inc_4n84) );
  INV_X4 vscale_core_DW01_inc_4_U284 ( .A(pipeline_csr_instret_full[29]), .ZN(vscale_core_DW01_inc_4n81) );
  INV_X4 vscale_core_DW01_inc_4_U285 ( .A(pipeline_csr_instret_full[30]), .ZN(vscale_core_DW01_inc_4n77) );
  INV_X4 vscale_core_DW01_inc_4_U286 ( .A(pipeline_csr_instret_full[31]), .ZN(vscale_core_DW01_inc_4n74) );
  INV_X4 vscale_core_DW01_inc_4_U287 ( .A(vscale_core_DW01_inc_4n68), .ZN(vscale_core_DW01_inc_4n67) );
  INV_X4 vscale_core_DW01_inc_4_U288 ( .A(pipeline_csr_instret_full[32]), .ZN(vscale_core_DW01_inc_4n66) );
  INV_X4 vscale_core_DW01_inc_4_U289 ( .A(pipeline_csr_instret_full[33]), .ZN(vscale_core_DW01_inc_4n63) );
  INV_X4 vscale_core_DW01_inc_4_U290 ( .A(vscale_core_DW01_inc_4n61), .ZN(vscale_core_DW01_inc_4n60) );
  INV_X4 vscale_core_DW01_inc_4_U291 ( .A(pipeline_csr_instret_full[34]), .ZN(vscale_core_DW01_inc_4n58) );
  INV_X4 vscale_core_DW01_inc_4_U292 ( .A(pipeline_csr_instret_full[35]), .ZN(vscale_core_DW01_inc_4n54) );
  INV_X4 vscale_core_DW01_inc_4_U293 ( .A(vscale_core_DW01_inc_4n50), .ZN(vscale_core_DW01_inc_4n49) );
  INV_X4 vscale_core_DW01_inc_4_U294 ( .A(pipeline_csr_instret_full[36]), .ZN(vscale_core_DW01_inc_4n48) );
  INV_X4 vscale_core_DW01_inc_4_U295 ( .A(pipeline_csr_instret_full[37]), .ZN(vscale_core_DW01_inc_4n44) );
  INV_X4 vscale_core_DW01_inc_4_U296 ( .A(vscale_core_DW01_inc_4n42), .ZN(vscale_core_DW01_inc_4n41) );
  INV_X4 vscale_core_DW01_inc_4_U297 ( .A(pipeline_csr_instret_full[38]), .ZN(vscale_core_DW01_inc_4n39) );
  INV_X4 vscale_core_DW01_inc_4_U298 ( .A(pipeline_csr_instret_full[39]), .ZN(vscale_core_DW01_inc_4n35) );
  INV_X4 vscale_core_DW01_inc_4_U299 ( .A(vscale_core_DW01_inc_4n31), .ZN(vscale_core_DW01_inc_4n30) );
  INV_X4 vscale_core_DW01_inc_4_U300 ( .A(n10618), .ZN(vscale_core_DW01_inc_4n28) );
  INV_X4 vscale_core_DW01_inc_4_U301 ( .A(pipeline_csr_instret_full[41]), .ZN(vscale_core_DW01_inc_4n25) );
  INV_X4 vscale_core_DW01_inc_4_U302 ( .A(pipeline_csr_instret_full[1]), .ZN(vscale_core_DW01_inc_4n203) );
  INV_X4 vscale_core_DW01_inc_4_U303 ( .A(vscale_core_DW01_inc_4n201), .ZN(vscale_core_DW01_inc_4n200) );
  INV_X4 vscale_core_DW01_inc_4_U304 ( .A(pipeline_csr_instret_full[2]), .ZN(vscale_core_DW01_inc_4n199) );
  INV_X4 vscale_core_DW01_inc_4_U305 ( .A(pipeline_csr_instret_full[3]), .ZN(vscale_core_DW01_inc_4n196) );
  INV_X4 vscale_core_DW01_inc_4_U306 ( .A(vscale_core_DW01_inc_4n193), .ZN(vscale_core_DW01_inc_4n192) );
  INV_X4 vscale_core_DW01_inc_4_U307 ( .A(pipeline_csr_instret_full[4]), .ZN(vscale_core_DW01_inc_4n191) );
  INV_X4 vscale_core_DW01_inc_4_U308 ( .A(pipeline_csr_instret_full[5]), .ZN(vscale_core_DW01_inc_4n187) );
  INV_X4 vscale_core_DW01_inc_4_U309 ( .A(pipeline_csr_instret_full[6]), .ZN(vscale_core_DW01_inc_4n183) );
  INV_X4 vscale_core_DW01_inc_4_U310 ( .A(pipeline_csr_instret_full[7]), .ZN(vscale_core_DW01_inc_4n180) );
  INV_X4 vscale_core_DW01_inc_4_U311 ( .A(vscale_core_DW01_inc_4n176), .ZN(vscale_core_DW01_inc_4n175) );
  INV_X4 vscale_core_DW01_inc_4_U312 ( .A(pipeline_csr_instret_full[8]), .ZN(vscale_core_DW01_inc_4n174) );
  INV_X4 vscale_core_DW01_inc_4_U313 ( .A(pipeline_csr_instret_full[9]), .ZN(vscale_core_DW01_inc_4n171) );
  INV_X4 vscale_core_DW01_inc_4_U314 ( .A(vscale_core_DW01_inc_4n169), .ZN(vscale_core_DW01_inc_4n168) );
  INV_X4 vscale_core_DW01_inc_4_U315 ( .A(pipeline_csr_instret_full[10]), .ZN(vscale_core_DW01_inc_4n166) );
  INV_X4 vscale_core_DW01_inc_4_U316 ( .A(pipeline_csr_instret_full[11]), .ZN(vscale_core_DW01_inc_4n162) );
  INV_X4 vscale_core_DW01_inc_4_U317 ( .A(vscale_core_DW01_inc_4n158), .ZN(vscale_core_DW01_inc_4n157) );
  INV_X4 vscale_core_DW01_inc_4_U318 ( .A(pipeline_csr_instret_full[12]), .ZN(vscale_core_DW01_inc_4n156) );
  INV_X4 vscale_core_DW01_inc_4_U319 ( .A(pipeline_csr_instret_full[13]), .ZN(vscale_core_DW01_inc_4n152) );
  INV_X4 vscale_core_DW01_inc_4_U320 ( .A(vscale_core_DW01_inc_4n150), .ZN(vscale_core_DW01_inc_4n149) );
  INV_X4 vscale_core_DW01_inc_4_U321 ( .A(pipeline_csr_instret_full[14]), .ZN(vscale_core_DW01_inc_4n147) );
  INV_X4 vscale_core_DW01_inc_4_U322 ( .A(pipeline_csr_instret_full[15]), .ZN(vscale_core_DW01_inc_4n143) );
  INV_X4 vscale_core_DW01_inc_4_U323 ( .A(vscale_core_DW01_inc_4n138), .ZN(vscale_core_DW01_inc_4n137) );
  INV_X4 vscale_core_DW01_inc_4_U324 ( .A(pipeline_csr_instret_full[16]), .ZN(vscale_core_DW01_inc_4n136) );
  INV_X4 vscale_core_DW01_inc_4_U325 ( .A(pipeline_csr_instret_full[17]), .ZN(vscale_core_DW01_inc_4n132) );
  INV_X4 vscale_core_DW01_inc_4_U326 ( .A(pipeline_csr_instret_full[18]), .ZN(vscale_core_DW01_inc_4n128) );
  INV_X4 vscale_core_DW01_inc_4_U327 ( .A(pipeline_csr_instret_full[19]), .ZN(vscale_core_DW01_inc_4n125) );
  INV_X4 vscale_core_DW01_inc_4_U328 ( .A(vscale_core_DW01_inc_4n122), .ZN(vscale_core_DW01_inc_4n121) );
  INV_X4 vscale_core_DW01_inc_4_U329 ( .A(vscale_core_DW01_inc_4n120), .ZN(vscale_core_DW01_inc_4n119) );
  INV_X4 vscale_core_DW01_inc_4_U330 ( .A(pipeline_csr_instret_full[20]), .ZN(vscale_core_DW01_inc_4n118) );
  INV_X4 vscale_core_DW01_inc_4_U331 ( .A(pipeline_csr_instret_full[21]), .ZN(vscale_core_DW01_inc_4n115) );
  INV_X4 vscale_core_DW01_inc_4_U332 ( .A(pipeline_csr_instret_full[22]), .ZN(vscale_core_DW01_inc_4n111) );
  INV_X4 vscale_core_DW01_inc_4_U333 ( .A(pipeline_csr_instret_full[23]), .ZN(vscale_core_DW01_inc_4n108) );
  INV_X4 vscale_core_DW01_inc_4_U334 ( .A(vscale_core_DW01_inc_4n103), .ZN(vscale_core_DW01_inc_4n102) );
  INV_X4 vscale_core_DW01_inc_4_U335 ( .A(pipeline_csr_instret_full[24]), .ZN(vscale_core_DW01_inc_4n101) );
;
  vscale_core_DW01_inc_5 pipeline_csr_add_315 

  XOR2_X2 vscale_core_DW01_inc_5_U1 ( .A(pipeline_csr_mtime_full[63]), .B(vscale_core_DW01_inc_5n1), .Z(pipeline_csr_N903) );
  HA_X1 vscale_core_DW01_inc_5_U2 ( .A(pipeline_csr_mtime_full[62]), .B(vscale_core_DW01_inc_5n2), .CO(vscale_core_DW01_inc_5n1), .S(pipeline_csr_N902) );
  HA_X1 vscale_core_DW01_inc_5_U3 ( .A(pipeline_csr_mtime_full[61]), .B(vscale_core_DW01_inc_5n3), .CO(vscale_core_DW01_inc_5n2), .S(pipeline_csr_N901) );
  HA_X1 vscale_core_DW01_inc_5_U4 ( .A(pipeline_csr_mtime_full[60]), .B(vscale_core_DW01_inc_5n4), .CO(vscale_core_DW01_inc_5n3), .S(pipeline_csr_N900) );
  HA_X1 vscale_core_DW01_inc_5_U5 ( .A(pipeline_csr_mtime_full[59]), .B(vscale_core_DW01_inc_5n5), .CO(vscale_core_DW01_inc_5n4), .S(pipeline_csr_N899) );
  HA_X1 vscale_core_DW01_inc_5_U6 ( .A(pipeline_csr_mtime_full[58]), .B(vscale_core_DW01_inc_5n6), .CO(vscale_core_DW01_inc_5n5), .S(pipeline_csr_N898) );
  HA_X1 vscale_core_DW01_inc_5_U7 ( .A(pipeline_csr_mtime_full[57]), .B(vscale_core_DW01_inc_5n7), .CO(vscale_core_DW01_inc_5n6), .S(pipeline_csr_N897) );
  HA_X1 vscale_core_DW01_inc_5_U8 ( .A(pipeline_csr_mtime_full[56]), .B(vscale_core_DW01_inc_5n8), .CO(vscale_core_DW01_inc_5n7), .S(pipeline_csr_N896) );
  HA_X1 vscale_core_DW01_inc_5_U9 ( .A(pipeline_csr_mtime_full[55]), .B(vscale_core_DW01_inc_5n9), .CO(vscale_core_DW01_inc_5n8), .S(pipeline_csr_N895) );
  HA_X1 vscale_core_DW01_inc_5_U10 ( .A(pipeline_csr_mtime_full[54]), .B(vscale_core_DW01_inc_5n10), .CO(vscale_core_DW01_inc_5n9), .S(pipeline_csr_N894) );
  HA_X1 vscale_core_DW01_inc_5_U11 ( .A(pipeline_csr_mtime_full[53]), .B(vscale_core_DW01_inc_5n11), .CO(vscale_core_DW01_inc_5n10), .S(pipeline_csr_N893) );
  HA_X1 vscale_core_DW01_inc_5_U12 ( .A(pipeline_csr_mtime_full[52]), .B(vscale_core_DW01_inc_5n12), .CO(vscale_core_DW01_inc_5n11), .S(pipeline_csr_N892) );
  HA_X1 vscale_core_DW01_inc_5_U13 ( .A(pipeline_csr_mtime_full[51]), .B(vscale_core_DW01_inc_5n13), .CO(vscale_core_DW01_inc_5n12), .S(pipeline_csr_N891) );
  HA_X1 vscale_core_DW01_inc_5_U14 ( .A(pipeline_csr_mtime_full[50]), .B(vscale_core_DW01_inc_5n14), .CO(vscale_core_DW01_inc_5n13), .S(pipeline_csr_N890) );
  HA_X1 vscale_core_DW01_inc_5_U15 ( .A(pipeline_csr_mtime_full[49]), .B(vscale_core_DW01_inc_5n15), .CO(vscale_core_DW01_inc_5n14), .S(pipeline_csr_N889) );
  HA_X1 vscale_core_DW01_inc_5_U16 ( .A(pipeline_csr_mtime_full[48]), .B(vscale_core_DW01_inc_5n16), .CO(vscale_core_DW01_inc_5n15), .S(pipeline_csr_N888) );
  HA_X1 vscale_core_DW01_inc_5_U17 ( .A(pipeline_csr_mtime_full[47]), .B(vscale_core_DW01_inc_5n17), .CO(vscale_core_DW01_inc_5n16), .S(pipeline_csr_N887) );
  HA_X1 vscale_core_DW01_inc_5_U18 ( .A(pipeline_csr_mtime_full[46]), .B(vscale_core_DW01_inc_5n18), .CO(vscale_core_DW01_inc_5n17), .S(pipeline_csr_N886) );
  HA_X1 vscale_core_DW01_inc_5_U19 ( .A(pipeline_csr_mtime_full[45]), .B(vscale_core_DW01_inc_5n19), .CO(vscale_core_DW01_inc_5n18), .S(pipeline_csr_N885) );
  HA_X1 vscale_core_DW01_inc_5_U20 ( .A(pipeline_csr_mtime_full[44]), .B(vscale_core_DW01_inc_5n20), .CO(vscale_core_DW01_inc_5n19), .S(pipeline_csr_N884) );
  HA_X1 vscale_core_DW01_inc_5_U21 ( .A(pipeline_csr_mtime_full[43]), .B(vscale_core_DW01_inc_5n21), .CO(vscale_core_DW01_inc_5n20), .S(pipeline_csr_N883) );
  HA_X1 vscale_core_DW01_inc_5_U22 ( .A(pipeline_csr_mtime_full[42]), .B(vscale_core_DW01_inc_5n22), .CO(vscale_core_DW01_inc_5n21), .S(pipeline_csr_N882) );
  XOR2_X2 vscale_core_DW01_inc_5_U23 ( .A(vscale_core_DW01_inc_5n25), .B(vscale_core_DW01_inc_5n26), .Z(pipeline_csr_N881) );
  NAND2_X2 vscale_core_DW01_inc_5_U25 ( .A1(vscale_core_DW01_inc_5n27), .A2(pipeline_csr_mtime_full[41]), .ZN(vscale_core_DW01_inc_5n23) );
  XOR2_X2 vscale_core_DW01_inc_5_U28 ( .A(vscale_core_DW01_inc_5n28), .B(vscale_core_DW01_inc_5n29), .Z(pipeline_csr_N880) );
  NAND2_X2 vscale_core_DW01_inc_5_U29 ( .A1(vscale_core_DW01_inc_5n67), .A2(vscale_core_DW01_inc_5n27), .ZN(vscale_core_DW01_inc_5n26) );
  XNOR2_X2 vscale_core_DW01_inc_5_U32 ( .A(vscale_core_DW01_inc_5n36), .B(vscale_core_DW01_inc_5n35), .ZN(pipeline_csr_N879) );
  NAND2_X2 vscale_core_DW01_inc_5_U33 ( .A1(vscale_core_DW01_inc_5n67), .A2(vscale_core_DW01_inc_5n30), .ZN(vscale_core_DW01_inc_5n29) );
  NAND2_X2 vscale_core_DW01_inc_5_U35 ( .A1(vscale_core_DW01_inc_5n51), .A2(vscale_core_DW01_inc_5n32), .ZN(vscale_core_DW01_inc_5n31) );
  NAND2_X2 vscale_core_DW01_inc_5_U37 ( .A1(pipeline_csr_mtime_full[38]), .A2(pipeline_csr_mtime_full[39]), .ZN(vscale_core_DW01_inc_5n33) );
  XOR2_X2 vscale_core_DW01_inc_5_U40 ( .A(vscale_core_DW01_inc_5n39), .B(vscale_core_DW01_inc_5n40), .Z(pipeline_csr_N878) );
  XNOR2_X2 vscale_core_DW01_inc_5_U45 ( .A(vscale_core_DW01_inc_5n45), .B(vscale_core_DW01_inc_5n44), .ZN(pipeline_csr_N877) );
  NAND2_X2 vscale_core_DW01_inc_5_U46 ( .A1(vscale_core_DW01_inc_5n49), .A2(vscale_core_DW01_inc_5n41), .ZN(vscale_core_DW01_inc_5n40) );
  NAND2_X2 vscale_core_DW01_inc_5_U48 ( .A1(pipeline_csr_mtime_full[36]), .A2(pipeline_csr_mtime_full[37]), .ZN(vscale_core_DW01_inc_5n42) );
  XNOR2_X2 vscale_core_DW01_inc_5_U51 ( .A(vscale_core_DW01_inc_5n49), .B(vscale_core_DW01_inc_5n48), .ZN(pipeline_csr_N876) );
  XNOR2_X2 vscale_core_DW01_inc_5_U56 ( .A(vscale_core_DW01_inc_5n55), .B(vscale_core_DW01_inc_5n54), .ZN(pipeline_csr_N875) );
  NAND2_X2 vscale_core_DW01_inc_5_U58 ( .A1(vscale_core_DW01_inc_5n67), .A2(vscale_core_DW01_inc_5n51), .ZN(vscale_core_DW01_inc_5n50) );
  NAND2_X2 vscale_core_DW01_inc_5_U60 ( .A1(pipeline_csr_mtime_full[34]), .A2(pipeline_csr_mtime_full[35]), .ZN(vscale_core_DW01_inc_5n52) );
  XOR2_X2 vscale_core_DW01_inc_5_U63 ( .A(vscale_core_DW01_inc_5n58), .B(vscale_core_DW01_inc_5n59), .Z(pipeline_csr_N874) );
  XOR2_X2 vscale_core_DW01_inc_5_U68 ( .A(vscale_core_DW01_inc_5n63), .B(vscale_core_DW01_inc_5n64), .Z(pipeline_csr_N873) );
  NAND2_X2 vscale_core_DW01_inc_5_U69 ( .A1(vscale_core_DW01_inc_5n67), .A2(vscale_core_DW01_inc_5n60), .ZN(vscale_core_DW01_inc_5n59) );
  NAND2_X2 vscale_core_DW01_inc_5_U71 ( .A1(pipeline_csr_mtime_full[32]), .A2(pipeline_csr_mtime_full[33]), .ZN(vscale_core_DW01_inc_5n61) );
  XNOR2_X2 vscale_core_DW01_inc_5_U74 ( .A(vscale_core_DW01_inc_5n67), .B(vscale_core_DW01_inc_5n66), .ZN(pipeline_csr_N872) );
  NAND2_X2 vscale_core_DW01_inc_5_U75 ( .A1(vscale_core_DW01_inc_5n67), .A2(pipeline_csr_mtime_full[32]), .ZN(vscale_core_DW01_inc_5n64) );
  XOR2_X2 vscale_core_DW01_inc_5_U78 ( .A(vscale_core_DW01_inc_5n74), .B(vscale_core_DW01_inc_5n75), .Z(pipeline_csr_N871) );
  NAND2_X2 vscale_core_DW01_inc_5_U80 ( .A1(vscale_core_DW01_inc_5n69), .A2(vscale_core_DW01_inc_5n138), .ZN(vscale_core_DW01_inc_5n68) );
  NAND2_X2 vscale_core_DW01_inc_5_U82 ( .A1(vscale_core_DW01_inc_5n88), .A2(vscale_core_DW01_inc_5n71), .ZN(vscale_core_DW01_inc_5n70) );
  NAND2_X2 vscale_core_DW01_inc_5_U84 ( .A1(pipeline_csr_mtime_full[30]), .A2(pipeline_csr_mtime_full[31]), .ZN(vscale_core_DW01_inc_5n72) );
  XNOR2_X2 vscale_core_DW01_inc_5_U87 ( .A(vscale_core_DW01_inc_5n78), .B(vscale_core_DW01_inc_5n77), .ZN(pipeline_csr_N870) );
  NAND2_X2 vscale_core_DW01_inc_5_U88 ( .A1(vscale_core_DW01_inc_5n78), .A2(pipeline_csr_mtime_full[30]), .ZN(vscale_core_DW01_inc_5n75) );
  XOR2_X2 vscale_core_DW01_inc_5_U91 ( .A(vscale_core_DW01_inc_5n81), .B(vscale_core_DW01_inc_5n82), .Z(pipeline_csr_N869) );
  NAND2_X2 vscale_core_DW01_inc_5_U93 ( .A1(pipeline_csr_mtime_full[28]), .A2(pipeline_csr_mtime_full[29]), .ZN(vscale_core_DW01_inc_5n79) );
  XOR2_X2 vscale_core_DW01_inc_5_U96 ( .A(vscale_core_DW01_inc_5n84), .B(vscale_core_DW01_inc_5n85), .Z(pipeline_csr_N868) );
  NAND2_X2 vscale_core_DW01_inc_5_U97 ( .A1(vscale_core_DW01_inc_5n86), .A2(pipeline_csr_mtime_full[28]), .ZN(vscale_core_DW01_inc_5n82) );
  XOR2_X2 vscale_core_DW01_inc_5_U100 ( .A(vscale_core_DW01_inc_5n91), .B(vscale_core_DW01_inc_5n92), .Z(pipeline_csr_N867) );
  NAND2_X2 vscale_core_DW01_inc_5_U105 ( .A1(pipeline_csr_mtime_full[26]), .A2(pipeline_csr_mtime_full[27]), .ZN(vscale_core_DW01_inc_5n89) );
  XNOR2_X2 vscale_core_DW01_inc_5_U108 ( .A(vscale_core_DW01_inc_5n95), .B(vscale_core_DW01_inc_5n94), .ZN(pipeline_csr_N866) );
  NAND2_X2 vscale_core_DW01_inc_5_U109 ( .A1(vscale_core_DW01_inc_5n95), .A2(pipeline_csr_mtime_full[26]), .ZN(vscale_core_DW01_inc_5n92) );
  XOR2_X2 vscale_core_DW01_inc_5_U112 ( .A(vscale_core_DW01_inc_5n98), .B(vscale_core_DW01_inc_5n99), .Z(pipeline_csr_N865) );
  NAND2_X2 vscale_core_DW01_inc_5_U114 ( .A1(pipeline_csr_mtime_full[24]), .A2(pipeline_csr_mtime_full[25]), .ZN(vscale_core_DW01_inc_5n96) );
  XOR2_X2 vscale_core_DW01_inc_5_U117 ( .A(vscale_core_DW01_inc_5n101), .B(vscale_core_DW01_inc_5n102), .Z(pipeline_csr_N864) );
  NAND2_X2 vscale_core_DW01_inc_5_U118 ( .A1(vscale_core_DW01_inc_5n103), .A2(pipeline_csr_mtime_full[24]), .ZN(vscale_core_DW01_inc_5n99) );
  XOR2_X2 vscale_core_DW01_inc_5_U121 ( .A(vscale_core_DW01_inc_5n108), .B(vscale_core_DW01_inc_5n109), .Z(pipeline_csr_N863) );
  NAND2_X2 vscale_core_DW01_inc_5_U124 ( .A1(vscale_core_DW01_inc_5n122), .A2(vscale_core_DW01_inc_5n105), .ZN(vscale_core_DW01_inc_5n104) );
  NAND2_X2 vscale_core_DW01_inc_5_U126 ( .A1(pipeline_csr_mtime_full[22]), .A2(pipeline_csr_mtime_full[23]), .ZN(vscale_core_DW01_inc_5n106) );
  XNOR2_X2 vscale_core_DW01_inc_5_U129 ( .A(vscale_core_DW01_inc_5n112), .B(vscale_core_DW01_inc_5n111), .ZN(pipeline_csr_N862) );
  NAND2_X2 vscale_core_DW01_inc_5_U130 ( .A1(vscale_core_DW01_inc_5n112), .A2(pipeline_csr_mtime_full[22]), .ZN(vscale_core_DW01_inc_5n109) );
  XOR2_X2 vscale_core_DW01_inc_5_U133 ( .A(vscale_core_DW01_inc_5n115), .B(vscale_core_DW01_inc_5n116), .Z(pipeline_csr_N861) );
  NAND2_X2 vscale_core_DW01_inc_5_U135 ( .A1(pipeline_csr_mtime_full[20]), .A2(pipeline_csr_mtime_full[21]), .ZN(vscale_core_DW01_inc_5n113) );
  XOR2_X2 vscale_core_DW01_inc_5_U138 ( .A(vscale_core_DW01_inc_5n118), .B(vscale_core_DW01_inc_5n119), .Z(pipeline_csr_N860) );
  NAND2_X2 vscale_core_DW01_inc_5_U139 ( .A1(vscale_core_DW01_inc_5n120), .A2(pipeline_csr_mtime_full[20]), .ZN(vscale_core_DW01_inc_5n116) );
  XOR2_X2 vscale_core_DW01_inc_5_U142 ( .A(vscale_core_DW01_inc_5n125), .B(vscale_core_DW01_inc_5n126), .Z(pipeline_csr_N859) );
  NAND2_X2 vscale_core_DW01_inc_5_U147 ( .A1(pipeline_csr_mtime_full[18]), .A2(pipeline_csr_mtime_full[19]), .ZN(vscale_core_DW01_inc_5n123) );
  XNOR2_X2 vscale_core_DW01_inc_5_U150 ( .A(vscale_core_DW01_inc_5n129), .B(vscale_core_DW01_inc_5n128), .ZN(pipeline_csr_N858) );
  NAND2_X2 vscale_core_DW01_inc_5_U151 ( .A1(vscale_core_DW01_inc_5n129), .A2(pipeline_csr_mtime_full[18]), .ZN(vscale_core_DW01_inc_5n126) );
  XNOR2_X2 vscale_core_DW01_inc_5_U154 ( .A(vscale_core_DW01_inc_5n133), .B(vscale_core_DW01_inc_5n132), .ZN(pipeline_csr_N857) );
  NAND2_X2 vscale_core_DW01_inc_5_U156 ( .A1(pipeline_csr_mtime_full[16]), .A2(pipeline_csr_mtime_full[17]), .ZN(vscale_core_DW01_inc_5n130) );
  XOR2_X2 vscale_core_DW01_inc_5_U159 ( .A(vscale_core_DW01_inc_5n136), .B(vscale_core_DW01_inc_5n137), .Z(pipeline_csr_N856) );
  XNOR2_X2 vscale_core_DW01_inc_5_U164 ( .A(vscale_core_DW01_inc_5n144), .B(vscale_core_DW01_inc_5n143), .ZN(pipeline_csr_N855) );
  NAND2_X2 vscale_core_DW01_inc_5_U167 ( .A1(vscale_core_DW01_inc_5n159), .A2(vscale_core_DW01_inc_5n140), .ZN(vscale_core_DW01_inc_5n139) );
  NAND2_X2 vscale_core_DW01_inc_5_U169 ( .A1(pipeline_csr_mtime_full[14]), .A2(pipeline_csr_mtime_full[15]), .ZN(vscale_core_DW01_inc_5n141) );
  XOR2_X2 vscale_core_DW01_inc_5_U172 ( .A(vscale_core_DW01_inc_5n147), .B(vscale_core_DW01_inc_5n148), .Z(pipeline_csr_N854) );
  XNOR2_X2 vscale_core_DW01_inc_5_U177 ( .A(vscale_core_DW01_inc_5n153), .B(vscale_core_DW01_inc_5n152), .ZN(pipeline_csr_N853) );
  NAND2_X2 vscale_core_DW01_inc_5_U178 ( .A1(vscale_core_DW01_inc_5n157), .A2(vscale_core_DW01_inc_5n149), .ZN(vscale_core_DW01_inc_5n148) );
  NAND2_X2 vscale_core_DW01_inc_5_U180 ( .A1(pipeline_csr_mtime_full[12]), .A2(pipeline_csr_mtime_full[13]), .ZN(vscale_core_DW01_inc_5n150) );
  XNOR2_X2 vscale_core_DW01_inc_5_U183 ( .A(vscale_core_DW01_inc_5n157), .B(vscale_core_DW01_inc_5n156), .ZN(pipeline_csr_N852) );
  XNOR2_X2 vscale_core_DW01_inc_5_U188 ( .A(vscale_core_DW01_inc_5n163), .B(vscale_core_DW01_inc_5n162), .ZN(pipeline_csr_N851) );
  NAND2_X2 vscale_core_DW01_inc_5_U190 ( .A1(vscale_core_DW01_inc_5n175), .A2(vscale_core_DW01_inc_5n159), .ZN(vscale_core_DW01_inc_5n158) );
  NAND2_X2 vscale_core_DW01_inc_5_U192 ( .A1(pipeline_csr_mtime_full[10]), .A2(pipeline_csr_mtime_full[11]), .ZN(vscale_core_DW01_inc_5n160) );
  XOR2_X2 vscale_core_DW01_inc_5_U195 ( .A(vscale_core_DW01_inc_5n166), .B(vscale_core_DW01_inc_5n167), .Z(pipeline_csr_N850) );
  XOR2_X2 vscale_core_DW01_inc_5_U200 ( .A(vscale_core_DW01_inc_5n171), .B(vscale_core_DW01_inc_5n172), .Z(pipeline_csr_N849) );
  NAND2_X2 vscale_core_DW01_inc_5_U201 ( .A1(vscale_core_DW01_inc_5n175), .A2(vscale_core_DW01_inc_5n168), .ZN(vscale_core_DW01_inc_5n167) );
  NAND2_X2 vscale_core_DW01_inc_5_U203 ( .A1(pipeline_csr_mtime_full[8]), .A2(pipeline_csr_mtime_full[9]), .ZN(vscale_core_DW01_inc_5n169) );
  XNOR2_X2 vscale_core_DW01_inc_5_U206 ( .A(vscale_core_DW01_inc_5n175), .B(vscale_core_DW01_inc_5n174), .ZN(pipeline_csr_N848) );
  NAND2_X2 vscale_core_DW01_inc_5_U207 ( .A1(vscale_core_DW01_inc_5n175), .A2(pipeline_csr_mtime_full[8]), .ZN(vscale_core_DW01_inc_5n172) );
  XOR2_X2 vscale_core_DW01_inc_5_U210 ( .A(vscale_core_DW01_inc_5n180), .B(vscale_core_DW01_inc_5n181), .Z(pipeline_csr_N847) );
  NAND2_X2 vscale_core_DW01_inc_5_U212 ( .A1(vscale_core_DW01_inc_5n177), .A2(vscale_core_DW01_inc_5n193), .ZN(vscale_core_DW01_inc_5n176) );
  NAND2_X2 vscale_core_DW01_inc_5_U214 ( .A1(pipeline_csr_mtime_full[6]), .A2(pipeline_csr_mtime_full[7]), .ZN(vscale_core_DW01_inc_5n178) );
  XNOR2_X2 vscale_core_DW01_inc_5_U217 ( .A(vscale_core_DW01_inc_5n184), .B(vscale_core_DW01_inc_5n183), .ZN(pipeline_csr_N846) );
  NAND2_X2 vscale_core_DW01_inc_5_U218 ( .A1(vscale_core_DW01_inc_5n184), .A2(pipeline_csr_mtime_full[6]), .ZN(vscale_core_DW01_inc_5n181) );
  XNOR2_X2 vscale_core_DW01_inc_5_U221 ( .A(vscale_core_DW01_inc_5n188), .B(vscale_core_DW01_inc_5n187), .ZN(pipeline_csr_N845) );
  NAND2_X2 vscale_core_DW01_inc_5_U223 ( .A1(pipeline_csr_mtime_full[4]), .A2(pipeline_csr_mtime_full[5]), .ZN(vscale_core_DW01_inc_5n185) );
  XOR2_X2 vscale_core_DW01_inc_5_U226 ( .A(vscale_core_DW01_inc_5n191), .B(vscale_core_DW01_inc_5n192), .Z(pipeline_csr_N844) );
  XOR2_X2 vscale_core_DW01_inc_5_U231 ( .A(vscale_core_DW01_inc_5n196), .B(vscale_core_DW01_inc_5n197), .Z(pipeline_csr_N843) );
  NAND2_X2 vscale_core_DW01_inc_5_U234 ( .A1(pipeline_csr_mtime_full[2]), .A2(pipeline_csr_mtime_full[3]), .ZN(vscale_core_DW01_inc_5n194) );
  XNOR2_X2 vscale_core_DW01_inc_5_U237 ( .A(vscale_core_DW01_inc_5n200), .B(vscale_core_DW01_inc_5n199), .ZN(pipeline_csr_N842) );
  NAND2_X2 vscale_core_DW01_inc_5_U238 ( .A1(vscale_core_DW01_inc_5n200), .A2(pipeline_csr_mtime_full[2]), .ZN(vscale_core_DW01_inc_5n197) );
  XNOR2_X2 vscale_core_DW01_inc_5_U241 ( .A(vscale_core_DW01_inc_5n203), .B(pipeline_csr_mtime_full[0]), .ZN(pipeline_csr_N841) );
  NAND2_X2 vscale_core_DW01_inc_5_U243 ( .A1(pipeline_csr_mtime_full[1]), .A2(pipeline_csr_mtime_full[0]), .ZN(vscale_core_DW01_inc_5n201) );
  NOR2_X2 vscale_core_DW01_inc_5_U250 ( .A1(vscale_core_DW01_inc_5n104), .A2(vscale_core_DW01_inc_5n70), .ZN(vscale_core_DW01_inc_5n69) );
  NOR2_X2 vscale_core_DW01_inc_5_U251 ( .A1(vscale_core_DW01_inc_5n79), .A2(vscale_core_DW01_inc_5n72), .ZN(vscale_core_DW01_inc_5n71) );
  NOR2_X2 vscale_core_DW01_inc_5_U252 ( .A1(vscale_core_DW01_inc_5n31), .A2(vscale_core_DW01_inc_5n28), .ZN(vscale_core_DW01_inc_5n27) );
  NOR2_X2 vscale_core_DW01_inc_5_U253 ( .A1(vscale_core_DW01_inc_5n137), .A2(vscale_core_DW01_inc_5n104), .ZN(vscale_core_DW01_inc_5n103) );
  NOR2_X2 vscale_core_DW01_inc_5_U254 ( .A1(vscale_core_DW01_inc_5n137), .A2(vscale_core_DW01_inc_5n121), .ZN(vscale_core_DW01_inc_5n120) );
  NOR2_X2 vscale_core_DW01_inc_5_U255 ( .A1(vscale_core_DW01_inc_5n102), .A2(vscale_core_DW01_inc_5n87), .ZN(vscale_core_DW01_inc_5n86) );
  NOR2_X2 vscale_core_DW01_inc_5_U256 ( .A1(vscale_core_DW01_inc_5n119), .A2(vscale_core_DW01_inc_5n113), .ZN(vscale_core_DW01_inc_5n112) );
  NOR2_X2 vscale_core_DW01_inc_5_U257 ( .A1(vscale_core_DW01_inc_5n102), .A2(vscale_core_DW01_inc_5n96), .ZN(vscale_core_DW01_inc_5n95) );
  NOR2_X2 vscale_core_DW01_inc_5_U258 ( .A1(vscale_core_DW01_inc_5n85), .A2(vscale_core_DW01_inc_5n79), .ZN(vscale_core_DW01_inc_5n78) );
  NOR2_X2 vscale_core_DW01_inc_5_U259 ( .A1(vscale_core_DW01_inc_5n192), .A2(vscale_core_DW01_inc_5n185), .ZN(vscale_core_DW01_inc_5n184) );
  NOR2_X2 vscale_core_DW01_inc_5_U260 ( .A1(vscale_core_DW01_inc_5n137), .A2(vscale_core_DW01_inc_5n130), .ZN(vscale_core_DW01_inc_5n129) );
  NOR2_X2 vscale_core_DW01_inc_5_U261 ( .A1(vscale_core_DW01_inc_5n192), .A2(vscale_core_DW01_inc_5n191), .ZN(vscale_core_DW01_inc_5n188) );
  NOR2_X2 vscale_core_DW01_inc_5_U262 ( .A1(vscale_core_DW01_inc_5n158), .A2(vscale_core_DW01_inc_5n156), .ZN(vscale_core_DW01_inc_5n153) );
  NOR2_X2 vscale_core_DW01_inc_5_U263 ( .A1(vscale_core_DW01_inc_5n167), .A2(vscale_core_DW01_inc_5n166), .ZN(vscale_core_DW01_inc_5n163) );
  NOR2_X2 vscale_core_DW01_inc_5_U264 ( .A1(vscale_core_DW01_inc_5n137), .A2(vscale_core_DW01_inc_5n136), .ZN(vscale_core_DW01_inc_5n133) );
  NOR2_X2 vscale_core_DW01_inc_5_U265 ( .A1(vscale_core_DW01_inc_5n148), .A2(vscale_core_DW01_inc_5n147), .ZN(vscale_core_DW01_inc_5n144) );
  NOR2_X2 vscale_core_DW01_inc_5_U266 ( .A1(vscale_core_DW01_inc_5n50), .A2(vscale_core_DW01_inc_5n48), .ZN(vscale_core_DW01_inc_5n45) );
  NOR2_X2 vscale_core_DW01_inc_5_U267 ( .A1(vscale_core_DW01_inc_5n40), .A2(vscale_core_DW01_inc_5n39), .ZN(vscale_core_DW01_inc_5n36) );
  NOR2_X2 vscale_core_DW01_inc_5_U268 ( .A1(vscale_core_DW01_inc_5n59), .A2(vscale_core_DW01_inc_5n58), .ZN(vscale_core_DW01_inc_5n55) );
  NOR2_X2 vscale_core_DW01_inc_5_U269 ( .A1(vscale_core_DW01_inc_5n113), .A2(vscale_core_DW01_inc_5n106), .ZN(vscale_core_DW01_inc_5n105) );
  NOR2_X2 vscale_core_DW01_inc_5_U270 ( .A1(vscale_core_DW01_inc_5n42), .A2(vscale_core_DW01_inc_5n33), .ZN(vscale_core_DW01_inc_5n32) );
  NOR2_X2 vscale_core_DW01_inc_5_U271 ( .A1(vscale_core_DW01_inc_5n185), .A2(vscale_core_DW01_inc_5n178), .ZN(vscale_core_DW01_inc_5n177) );
  NOR2_X2 vscale_core_DW01_inc_5_U272 ( .A1(vscale_core_DW01_inc_5n68), .A2(vscale_core_DW01_inc_5n23), .ZN(vscale_core_DW01_inc_5n22) );
  NOR2_X2 vscale_core_DW01_inc_5_U273 ( .A1(vscale_core_DW01_inc_5n96), .A2(vscale_core_DW01_inc_5n89), .ZN(vscale_core_DW01_inc_5n88) );
  NOR2_X2 vscale_core_DW01_inc_5_U274 ( .A1(vscale_core_DW01_inc_5n130), .A2(vscale_core_DW01_inc_5n123), .ZN(vscale_core_DW01_inc_5n122) );
  NOR2_X2 vscale_core_DW01_inc_5_U275 ( .A1(vscale_core_DW01_inc_5n194), .A2(vscale_core_DW01_inc_5n201), .ZN(vscale_core_DW01_inc_5n193) );
  NOR2_X2 vscale_core_DW01_inc_5_U276 ( .A1(vscale_core_DW01_inc_5n139), .A2(vscale_core_DW01_inc_5n176), .ZN(vscale_core_DW01_inc_5n138) );
  NOR2_X2 vscale_core_DW01_inc_5_U277 ( .A1(vscale_core_DW01_inc_5n150), .A2(vscale_core_DW01_inc_5n141), .ZN(vscale_core_DW01_inc_5n140) );
  NOR2_X2 vscale_core_DW01_inc_5_U278 ( .A1(vscale_core_DW01_inc_5n169), .A2(vscale_core_DW01_inc_5n160), .ZN(vscale_core_DW01_inc_5n159) );
  NOR2_X2 vscale_core_DW01_inc_5_U279 ( .A1(vscale_core_DW01_inc_5n61), .A2(vscale_core_DW01_inc_5n52), .ZN(vscale_core_DW01_inc_5n51) );
  INV_X4 vscale_core_DW01_inc_5_U280 ( .A(pipeline_csr_mtime_full[25]), .ZN(vscale_core_DW01_inc_5n98) );
  INV_X4 vscale_core_DW01_inc_5_U281 ( .A(pipeline_csr_mtime_full[26]), .ZN(vscale_core_DW01_inc_5n94) );
  INV_X4 vscale_core_DW01_inc_5_U282 ( .A(pipeline_csr_mtime_full[27]), .ZN(vscale_core_DW01_inc_5n91) );
  INV_X4 vscale_core_DW01_inc_5_U283 ( .A(vscale_core_DW01_inc_5n88), .ZN(vscale_core_DW01_inc_5n87) );
  INV_X4 vscale_core_DW01_inc_5_U284 ( .A(vscale_core_DW01_inc_5n86), .ZN(vscale_core_DW01_inc_5n85) );
  INV_X4 vscale_core_DW01_inc_5_U285 ( .A(pipeline_csr_mtime_full[28]), .ZN(vscale_core_DW01_inc_5n84) );
  INV_X4 vscale_core_DW01_inc_5_U286 ( .A(pipeline_csr_mtime_full[29]), .ZN(vscale_core_DW01_inc_5n81) );
  INV_X4 vscale_core_DW01_inc_5_U287 ( .A(pipeline_csr_mtime_full[30]), .ZN(vscale_core_DW01_inc_5n77) );
  INV_X4 vscale_core_DW01_inc_5_U288 ( .A(pipeline_csr_mtime_full[31]), .ZN(vscale_core_DW01_inc_5n74) );
  INV_X4 vscale_core_DW01_inc_5_U289 ( .A(vscale_core_DW01_inc_5n68), .ZN(vscale_core_DW01_inc_5n67) );
  INV_X4 vscale_core_DW01_inc_5_U290 ( .A(pipeline_csr_mtime_full[32]), .ZN(vscale_core_DW01_inc_5n66) );
  INV_X4 vscale_core_DW01_inc_5_U291 ( .A(pipeline_csr_mtime_full[33]), .ZN(vscale_core_DW01_inc_5n63) );
  INV_X4 vscale_core_DW01_inc_5_U292 ( .A(vscale_core_DW01_inc_5n61), .ZN(vscale_core_DW01_inc_5n60) );
  INV_X4 vscale_core_DW01_inc_5_U293 ( .A(pipeline_csr_mtime_full[34]), .ZN(vscale_core_DW01_inc_5n58) );
  INV_X4 vscale_core_DW01_inc_5_U294 ( .A(pipeline_csr_mtime_full[35]), .ZN(vscale_core_DW01_inc_5n54) );
  INV_X4 vscale_core_DW01_inc_5_U295 ( .A(vscale_core_DW01_inc_5n50), .ZN(vscale_core_DW01_inc_5n49) );
  INV_X4 vscale_core_DW01_inc_5_U296 ( .A(pipeline_csr_mtime_full[36]), .ZN(vscale_core_DW01_inc_5n48) );
  INV_X4 vscale_core_DW01_inc_5_U297 ( .A(pipeline_csr_mtime_full[37]), .ZN(vscale_core_DW01_inc_5n44) );
  INV_X4 vscale_core_DW01_inc_5_U298 ( .A(vscale_core_DW01_inc_5n42), .ZN(vscale_core_DW01_inc_5n41) );
  INV_X4 vscale_core_DW01_inc_5_U299 ( .A(pipeline_csr_mtime_full[38]), .ZN(vscale_core_DW01_inc_5n39) );
  INV_X4 vscale_core_DW01_inc_5_U300 ( .A(pipeline_csr_mtime_full[39]), .ZN(vscale_core_DW01_inc_5n35) );
  INV_X4 vscale_core_DW01_inc_5_U301 ( .A(vscale_core_DW01_inc_5n31), .ZN(vscale_core_DW01_inc_5n30) );
  INV_X4 vscale_core_DW01_inc_5_U302 ( .A(pipeline_csr_mtime_full[40]), .ZN(vscale_core_DW01_inc_5n28) );
  INV_X4 vscale_core_DW01_inc_5_U303 ( .A(pipeline_csr_mtime_full[41]), .ZN(vscale_core_DW01_inc_5n25) );
  INV_X4 vscale_core_DW01_inc_5_U304 ( .A(pipeline_csr_mtime_full[1]), .ZN(vscale_core_DW01_inc_5n203) );
  INV_X4 vscale_core_DW01_inc_5_U305 ( .A(vscale_core_DW01_inc_5n201), .ZN(vscale_core_DW01_inc_5n200) );
  INV_X4 vscale_core_DW01_inc_5_U306 ( .A(pipeline_csr_mtime_full[2]), .ZN(vscale_core_DW01_inc_5n199) );
  INV_X4 vscale_core_DW01_inc_5_U307 ( .A(pipeline_csr_mtime_full[3]), .ZN(vscale_core_DW01_inc_5n196) );
  INV_X4 vscale_core_DW01_inc_5_U308 ( .A(vscale_core_DW01_inc_5n193), .ZN(vscale_core_DW01_inc_5n192) );
  INV_X4 vscale_core_DW01_inc_5_U309 ( .A(pipeline_csr_mtime_full[4]), .ZN(vscale_core_DW01_inc_5n191) );
  INV_X4 vscale_core_DW01_inc_5_U310 ( .A(pipeline_csr_mtime_full[5]), .ZN(vscale_core_DW01_inc_5n187) );
  INV_X4 vscale_core_DW01_inc_5_U311 ( .A(pipeline_csr_mtime_full[6]), .ZN(vscale_core_DW01_inc_5n183) );
  INV_X4 vscale_core_DW01_inc_5_U312 ( .A(pipeline_csr_mtime_full[7]), .ZN(vscale_core_DW01_inc_5n180) );
  INV_X4 vscale_core_DW01_inc_5_U313 ( .A(vscale_core_DW01_inc_5n176), .ZN(vscale_core_DW01_inc_5n175) );
  INV_X4 vscale_core_DW01_inc_5_U314 ( .A(pipeline_csr_mtime_full[8]), .ZN(vscale_core_DW01_inc_5n174) );
  INV_X4 vscale_core_DW01_inc_5_U315 ( .A(pipeline_csr_mtime_full[9]), .ZN(vscale_core_DW01_inc_5n171) );
  INV_X4 vscale_core_DW01_inc_5_U316 ( .A(vscale_core_DW01_inc_5n169), .ZN(vscale_core_DW01_inc_5n168) );
  INV_X4 vscale_core_DW01_inc_5_U317 ( .A(pipeline_csr_mtime_full[10]), .ZN(vscale_core_DW01_inc_5n166) );
  INV_X4 vscale_core_DW01_inc_5_U318 ( .A(pipeline_csr_mtime_full[11]), .ZN(vscale_core_DW01_inc_5n162) );
  INV_X4 vscale_core_DW01_inc_5_U319 ( .A(vscale_core_DW01_inc_5n158), .ZN(vscale_core_DW01_inc_5n157) );
  INV_X4 vscale_core_DW01_inc_5_U320 ( .A(pipeline_csr_mtime_full[12]), .ZN(vscale_core_DW01_inc_5n156) );
  INV_X4 vscale_core_DW01_inc_5_U321 ( .A(pipeline_csr_mtime_full[13]), .ZN(vscale_core_DW01_inc_5n152) );
  INV_X4 vscale_core_DW01_inc_5_U322 ( .A(vscale_core_DW01_inc_5n150), .ZN(vscale_core_DW01_inc_5n149) );
  INV_X4 vscale_core_DW01_inc_5_U323 ( .A(pipeline_csr_mtime_full[14]), .ZN(vscale_core_DW01_inc_5n147) );
  INV_X4 vscale_core_DW01_inc_5_U324 ( .A(pipeline_csr_mtime_full[15]), .ZN(vscale_core_DW01_inc_5n143) );
  INV_X4 vscale_core_DW01_inc_5_U325 ( .A(vscale_core_DW01_inc_5n138), .ZN(vscale_core_DW01_inc_5n137) );
  INV_X4 vscale_core_DW01_inc_5_U326 ( .A(pipeline_csr_mtime_full[16]), .ZN(vscale_core_DW01_inc_5n136) );
  INV_X4 vscale_core_DW01_inc_5_U327 ( .A(pipeline_csr_mtime_full[17]), .ZN(vscale_core_DW01_inc_5n132) );
  INV_X4 vscale_core_DW01_inc_5_U328 ( .A(pipeline_csr_mtime_full[18]), .ZN(vscale_core_DW01_inc_5n128) );
  INV_X4 vscale_core_DW01_inc_5_U329 ( .A(pipeline_csr_mtime_full[19]), .ZN(vscale_core_DW01_inc_5n125) );
  INV_X4 vscale_core_DW01_inc_5_U330 ( .A(vscale_core_DW01_inc_5n122), .ZN(vscale_core_DW01_inc_5n121) );
  INV_X4 vscale_core_DW01_inc_5_U331 ( .A(vscale_core_DW01_inc_5n120), .ZN(vscale_core_DW01_inc_5n119) );
  INV_X4 vscale_core_DW01_inc_5_U332 ( .A(pipeline_csr_mtime_full[20]), .ZN(vscale_core_DW01_inc_5n118) );
  INV_X4 vscale_core_DW01_inc_5_U333 ( .A(pipeline_csr_mtime_full[21]), .ZN(vscale_core_DW01_inc_5n115) );
  INV_X4 vscale_core_DW01_inc_5_U334 ( .A(pipeline_csr_mtime_full[22]), .ZN(vscale_core_DW01_inc_5n111) );
  INV_X4 vscale_core_DW01_inc_5_U335 ( .A(pipeline_csr_mtime_full[23]), .ZN(vscale_core_DW01_inc_5n108) );
  INV_X4 vscale_core_DW01_inc_5_U336 ( .A(vscale_core_DW01_inc_5n103), .ZN(vscale_core_DW01_inc_5n102) );
  INV_X4 vscale_core_DW01_inc_5_U337 ( .A(pipeline_csr_mtime_full[24]), .ZN(vscale_core_DW01_inc_5n101) );
  INV_X4 vscale_core_DW01_inc_5_U338 ( .A(pipeline_csr_mtime_full[0]), .ZN(pipeline_csr_N840) );
;
  vscale_core_DW01_inc_6 pipeline_csr_add_312 

  XOR2_X2 vscale_core_DW01_inc_6_U1 ( .A(pipeline_csr_time_full[63]), .B(vscale_core_DW01_inc_6n1), .Z(pipeline_csr_N775) );
  HA_X1 vscale_core_DW01_inc_6_U2 ( .A(pipeline_csr_time_full[62]), .B(vscale_core_DW01_inc_6n2), .CO(vscale_core_DW01_inc_6n1), .S(pipeline_csr_N774) );
  HA_X1 vscale_core_DW01_inc_6_U3 ( .A(pipeline_csr_time_full[61]), .B(vscale_core_DW01_inc_6n3), .CO(vscale_core_DW01_inc_6n2), .S(pipeline_csr_N773) );
  HA_X1 vscale_core_DW01_inc_6_U4 ( .A(pipeline_csr_time_full[60]), .B(vscale_core_DW01_inc_6n4), .CO(vscale_core_DW01_inc_6n3), .S(pipeline_csr_N772) );
  HA_X1 vscale_core_DW01_inc_6_U5 ( .A(pipeline_csr_time_full[59]), .B(vscale_core_DW01_inc_6n5), .CO(vscale_core_DW01_inc_6n4), .S(pipeline_csr_N771) );
  HA_X1 vscale_core_DW01_inc_6_U6 ( .A(pipeline_csr_time_full[58]), .B(vscale_core_DW01_inc_6n6), .CO(vscale_core_DW01_inc_6n5), .S(pipeline_csr_N770) );
  HA_X1 vscale_core_DW01_inc_6_U7 ( .A(pipeline_csr_time_full[57]), .B(vscale_core_DW01_inc_6n7), .CO(vscale_core_DW01_inc_6n6), .S(pipeline_csr_N769) );
  HA_X1 vscale_core_DW01_inc_6_U8 ( .A(pipeline_csr_time_full[56]), .B(vscale_core_DW01_inc_6n8), .CO(vscale_core_DW01_inc_6n7), .S(pipeline_csr_N768) );
  HA_X1 vscale_core_DW01_inc_6_U9 ( .A(pipeline_csr_time_full[55]), .B(vscale_core_DW01_inc_6n9), .CO(vscale_core_DW01_inc_6n8), .S(pipeline_csr_N767) );
  HA_X1 vscale_core_DW01_inc_6_U10 ( .A(pipeline_csr_time_full[54]), .B(vscale_core_DW01_inc_6n10), .CO(vscale_core_DW01_inc_6n9), .S(pipeline_csr_N766) );
  HA_X1 vscale_core_DW01_inc_6_U11 ( .A(pipeline_csr_time_full[53]), .B(vscale_core_DW01_inc_6n11), .CO(vscale_core_DW01_inc_6n10), .S(pipeline_csr_N765) );
  HA_X1 vscale_core_DW01_inc_6_U12 ( .A(pipeline_csr_time_full[52]), .B(vscale_core_DW01_inc_6n12), .CO(vscale_core_DW01_inc_6n11), .S(pipeline_csr_N764) );
  HA_X1 vscale_core_DW01_inc_6_U13 ( .A(pipeline_csr_time_full[51]), .B(vscale_core_DW01_inc_6n13), .CO(vscale_core_DW01_inc_6n12), .S(pipeline_csr_N763) );
  HA_X1 vscale_core_DW01_inc_6_U14 ( .A(pipeline_csr_time_full[50]), .B(vscale_core_DW01_inc_6n14), .CO(vscale_core_DW01_inc_6n13), .S(pipeline_csr_N762) );
  HA_X1 vscale_core_DW01_inc_6_U15 ( .A(pipeline_csr_time_full[49]), .B(vscale_core_DW01_inc_6n15), .CO(vscale_core_DW01_inc_6n14), .S(pipeline_csr_N761) );
  HA_X1 vscale_core_DW01_inc_6_U16 ( .A(pipeline_csr_time_full[48]), .B(vscale_core_DW01_inc_6n16), .CO(vscale_core_DW01_inc_6n15), .S(pipeline_csr_N760) );
  HA_X1 vscale_core_DW01_inc_6_U17 ( .A(pipeline_csr_time_full[47]), .B(vscale_core_DW01_inc_6n17), .CO(vscale_core_DW01_inc_6n16), .S(pipeline_csr_N759) );
  HA_X1 vscale_core_DW01_inc_6_U18 ( .A(pipeline_csr_time_full[46]), .B(vscale_core_DW01_inc_6n18), .CO(vscale_core_DW01_inc_6n17), .S(pipeline_csr_N758) );
  HA_X1 vscale_core_DW01_inc_6_U19 ( .A(pipeline_csr_time_full[45]), .B(vscale_core_DW01_inc_6n19), .CO(vscale_core_DW01_inc_6n18), .S(pipeline_csr_N757) );
  HA_X1 vscale_core_DW01_inc_6_U20 ( .A(pipeline_csr_time_full[44]), .B(vscale_core_DW01_inc_6n20), .CO(vscale_core_DW01_inc_6n19), .S(pipeline_csr_N756) );
  HA_X1 vscale_core_DW01_inc_6_U21 ( .A(pipeline_csr_time_full[43]), .B(vscale_core_DW01_inc_6n21), .CO(vscale_core_DW01_inc_6n20), .S(pipeline_csr_N755) );
  HA_X1 vscale_core_DW01_inc_6_U22 ( .A(pipeline_csr_time_full[42]), .B(vscale_core_DW01_inc_6n22), .CO(vscale_core_DW01_inc_6n21), .S(pipeline_csr_N754) );
  HA_X1 vscale_core_DW01_inc_6_U23 ( .A(pipeline_csr_time_full[41]), .B(vscale_core_DW01_inc_6n23), .CO(vscale_core_DW01_inc_6n22), .S(pipeline_csr_N753) );
  XOR2_X2 vscale_core_DW01_inc_6_U24 ( .A(vscale_core_DW01_inc_6n26), .B(vscale_core_DW01_inc_6n27), .Z(pipeline_csr_N752) );
  NAND2_X2 vscale_core_DW01_inc_6_U26 ( .A1(vscale_core_DW01_inc_6n28), .A2(pipeline_csr_time_full[40]), .ZN(vscale_core_DW01_inc_6n24) );
  XOR2_X2 vscale_core_DW01_inc_6_U29 ( .A(vscale_core_DW01_inc_6n29), .B(vscale_core_DW01_inc_6n30), .Z(pipeline_csr_N751) );
  NAND2_X2 vscale_core_DW01_inc_6_U30 ( .A1(vscale_core_DW01_inc_6n62), .A2(vscale_core_DW01_inc_6n28), .ZN(vscale_core_DW01_inc_6n27) );
  XOR2_X2 vscale_core_DW01_inc_6_U33 ( .A(vscale_core_DW01_inc_6n34), .B(vscale_core_DW01_inc_6n35), .Z(pipeline_csr_N750) );
  NAND2_X2 vscale_core_DW01_inc_6_U34 ( .A1(vscale_core_DW01_inc_6n62), .A2(vscale_core_DW01_inc_6n31), .ZN(vscale_core_DW01_inc_6n30) );
  NAND2_X2 vscale_core_DW01_inc_6_U36 ( .A1(vscale_core_DW01_inc_6n46), .A2(vscale_core_DW01_inc_6n33), .ZN(vscale_core_DW01_inc_6n32) );
  XNOR2_X2 vscale_core_DW01_inc_6_U39 ( .A(vscale_core_DW01_inc_6n40), .B(vscale_core_DW01_inc_6n39), .ZN(pipeline_csr_N749) );
  NAND2_X2 vscale_core_DW01_inc_6_U40 ( .A1(vscale_core_DW01_inc_6n44), .A2(vscale_core_DW01_inc_6n36), .ZN(vscale_core_DW01_inc_6n35) );
  NAND2_X2 vscale_core_DW01_inc_6_U42 ( .A1(pipeline_csr_time_full[36]), .A2(pipeline_csr_time_full[37]), .ZN(vscale_core_DW01_inc_6n37) );
  XNOR2_X2 vscale_core_DW01_inc_6_U45 ( .A(vscale_core_DW01_inc_6n44), .B(vscale_core_DW01_inc_6n43), .ZN(pipeline_csr_N748) );
  XNOR2_X2 vscale_core_DW01_inc_6_U50 ( .A(vscale_core_DW01_inc_6n50), .B(vscale_core_DW01_inc_6n49), .ZN(pipeline_csr_N747) );
  NAND2_X2 vscale_core_DW01_inc_6_U52 ( .A1(vscale_core_DW01_inc_6n62), .A2(vscale_core_DW01_inc_6n46), .ZN(vscale_core_DW01_inc_6n45) );
  NAND2_X2 vscale_core_DW01_inc_6_U54 ( .A1(pipeline_csr_time_full[34]), .A2(pipeline_csr_time_full[35]), .ZN(vscale_core_DW01_inc_6n47) );
  XOR2_X2 vscale_core_DW01_inc_6_U57 ( .A(vscale_core_DW01_inc_6n53), .B(vscale_core_DW01_inc_6n54), .Z(pipeline_csr_N746) );
  XOR2_X2 vscale_core_DW01_inc_6_U62 ( .A(vscale_core_DW01_inc_6n58), .B(vscale_core_DW01_inc_6n59), .Z(pipeline_csr_N745) );
  NAND2_X2 vscale_core_DW01_inc_6_U63 ( .A1(vscale_core_DW01_inc_6n62), .A2(vscale_core_DW01_inc_6n55), .ZN(vscale_core_DW01_inc_6n54) );
  NAND2_X2 vscale_core_DW01_inc_6_U65 ( .A1(pipeline_csr_time_full[32]), .A2(pipeline_csr_time_full[33]), .ZN(vscale_core_DW01_inc_6n56) );
  XNOR2_X2 vscale_core_DW01_inc_6_U68 ( .A(vscale_core_DW01_inc_6n62), .B(vscale_core_DW01_inc_6n61), .ZN(pipeline_csr_N744) );
  NAND2_X2 vscale_core_DW01_inc_6_U69 ( .A1(vscale_core_DW01_inc_6n62), .A2(pipeline_csr_time_full[32]), .ZN(vscale_core_DW01_inc_6n59) );
  XOR2_X2 vscale_core_DW01_inc_6_U72 ( .A(vscale_core_DW01_inc_6n69), .B(vscale_core_DW01_inc_6n70), .Z(pipeline_csr_N743) );
  NAND2_X2 vscale_core_DW01_inc_6_U74 ( .A1(vscale_core_DW01_inc_6n64), .A2(vscale_core_DW01_inc_6n133), .ZN(vscale_core_DW01_inc_6n63) );
  NAND2_X2 vscale_core_DW01_inc_6_U76 ( .A1(vscale_core_DW01_inc_6n83), .A2(vscale_core_DW01_inc_6n66), .ZN(vscale_core_DW01_inc_6n65) );
  NAND2_X2 vscale_core_DW01_inc_6_U78 ( .A1(pipeline_csr_time_full[30]), .A2(pipeline_csr_time_full[31]), .ZN(vscale_core_DW01_inc_6n67) );
  XNOR2_X2 vscale_core_DW01_inc_6_U81 ( .A(vscale_core_DW01_inc_6n73), .B(vscale_core_DW01_inc_6n72), .ZN(pipeline_csr_N742) );
  NAND2_X2 vscale_core_DW01_inc_6_U82 ( .A1(vscale_core_DW01_inc_6n73), .A2(pipeline_csr_time_full[30]), .ZN(vscale_core_DW01_inc_6n70) );
  XOR2_X2 vscale_core_DW01_inc_6_U85 ( .A(vscale_core_DW01_inc_6n76), .B(vscale_core_DW01_inc_6n77), .Z(pipeline_csr_N741) );
  NAND2_X2 vscale_core_DW01_inc_6_U87 ( .A1(pipeline_csr_time_full[28]), .A2(pipeline_csr_time_full[29]), .ZN(vscale_core_DW01_inc_6n74) );
  XOR2_X2 vscale_core_DW01_inc_6_U90 ( .A(vscale_core_DW01_inc_6n79), .B(vscale_core_DW01_inc_6n80), .Z(pipeline_csr_N740) );
  NAND2_X2 vscale_core_DW01_inc_6_U91 ( .A1(vscale_core_DW01_inc_6n81), .A2(pipeline_csr_time_full[28]), .ZN(vscale_core_DW01_inc_6n77) );
  XOR2_X2 vscale_core_DW01_inc_6_U94 ( .A(vscale_core_DW01_inc_6n86), .B(vscale_core_DW01_inc_6n87), .Z(pipeline_csr_N739) );
  NAND2_X2 vscale_core_DW01_inc_6_U99 ( .A1(pipeline_csr_time_full[26]), .A2(pipeline_csr_time_full[27]), .ZN(vscale_core_DW01_inc_6n84) );
  XNOR2_X2 vscale_core_DW01_inc_6_U102 ( .A(vscale_core_DW01_inc_6n90), .B(vscale_core_DW01_inc_6n89), .ZN(pipeline_csr_N738) );
  NAND2_X2 vscale_core_DW01_inc_6_U103 ( .A1(vscale_core_DW01_inc_6n90), .A2(pipeline_csr_time_full[26]), .ZN(vscale_core_DW01_inc_6n87) );
  XOR2_X2 vscale_core_DW01_inc_6_U106 ( .A(vscale_core_DW01_inc_6n93), .B(vscale_core_DW01_inc_6n94), .Z(pipeline_csr_N737) );
  NAND2_X2 vscale_core_DW01_inc_6_U108 ( .A1(pipeline_csr_time_full[24]), .A2(pipeline_csr_time_full[25]), .ZN(vscale_core_DW01_inc_6n91) );
  XOR2_X2 vscale_core_DW01_inc_6_U111 ( .A(vscale_core_DW01_inc_6n96), .B(vscale_core_DW01_inc_6n97), .Z(pipeline_csr_N736) );
  NAND2_X2 vscale_core_DW01_inc_6_U112 ( .A1(vscale_core_DW01_inc_6n98), .A2(pipeline_csr_time_full[24]), .ZN(vscale_core_DW01_inc_6n94) );
  XOR2_X2 vscale_core_DW01_inc_6_U115 ( .A(vscale_core_DW01_inc_6n103), .B(vscale_core_DW01_inc_6n104), .Z(pipeline_csr_N735) );
  NAND2_X2 vscale_core_DW01_inc_6_U118 ( .A1(vscale_core_DW01_inc_6n117), .A2(vscale_core_DW01_inc_6n100), .ZN(vscale_core_DW01_inc_6n99) );
  NAND2_X2 vscale_core_DW01_inc_6_U120 ( .A1(pipeline_csr_time_full[22]), .A2(pipeline_csr_time_full[23]), .ZN(vscale_core_DW01_inc_6n101) );
  XNOR2_X2 vscale_core_DW01_inc_6_U123 ( .A(vscale_core_DW01_inc_6n107), .B(vscale_core_DW01_inc_6n106), .ZN(pipeline_csr_N734) );
  NAND2_X2 vscale_core_DW01_inc_6_U124 ( .A1(vscale_core_DW01_inc_6n107), .A2(pipeline_csr_time_full[22]), .ZN(vscale_core_DW01_inc_6n104) );
  XOR2_X2 vscale_core_DW01_inc_6_U127 ( .A(vscale_core_DW01_inc_6n110), .B(vscale_core_DW01_inc_6n111), .Z(pipeline_csr_N733) );
  NAND2_X2 vscale_core_DW01_inc_6_U129 ( .A1(pipeline_csr_time_full[20]), .A2(pipeline_csr_time_full[21]), .ZN(vscale_core_DW01_inc_6n108) );
  XOR2_X2 vscale_core_DW01_inc_6_U132 ( .A(vscale_core_DW01_inc_6n113), .B(vscale_core_DW01_inc_6n114), .Z(pipeline_csr_N732) );
  NAND2_X2 vscale_core_DW01_inc_6_U133 ( .A1(vscale_core_DW01_inc_6n115), .A2(pipeline_csr_time_full[20]), .ZN(vscale_core_DW01_inc_6n111) );
  XOR2_X2 vscale_core_DW01_inc_6_U136 ( .A(vscale_core_DW01_inc_6n120), .B(vscale_core_DW01_inc_6n121), .Z(pipeline_csr_N731) );
  NAND2_X2 vscale_core_DW01_inc_6_U141 ( .A1(pipeline_csr_time_full[18]), .A2(pipeline_csr_time_full[19]), .ZN(vscale_core_DW01_inc_6n118) );
  XNOR2_X2 vscale_core_DW01_inc_6_U144 ( .A(vscale_core_DW01_inc_6n124), .B(vscale_core_DW01_inc_6n123), .ZN(pipeline_csr_N730) );
  NAND2_X2 vscale_core_DW01_inc_6_U145 ( .A1(vscale_core_DW01_inc_6n124), .A2(pipeline_csr_time_full[18]), .ZN(vscale_core_DW01_inc_6n121) );
  XNOR2_X2 vscale_core_DW01_inc_6_U148 ( .A(vscale_core_DW01_inc_6n128), .B(vscale_core_DW01_inc_6n127), .ZN(pipeline_csr_N729) );
  NAND2_X2 vscale_core_DW01_inc_6_U150 ( .A1(pipeline_csr_time_full[16]), .A2(pipeline_csr_time_full[17]), .ZN(vscale_core_DW01_inc_6n125) );
  XOR2_X2 vscale_core_DW01_inc_6_U153 ( .A(vscale_core_DW01_inc_6n131), .B(vscale_core_DW01_inc_6n132), .Z(pipeline_csr_N728) );
  XNOR2_X2 vscale_core_DW01_inc_6_U158 ( .A(vscale_core_DW01_inc_6n139), .B(vscale_core_DW01_inc_6n138), .ZN(pipeline_csr_N727) );
  NAND2_X2 vscale_core_DW01_inc_6_U161 ( .A1(vscale_core_DW01_inc_6n154), .A2(vscale_core_DW01_inc_6n135), .ZN(vscale_core_DW01_inc_6n134) );
  NAND2_X2 vscale_core_DW01_inc_6_U163 ( .A1(pipeline_csr_time_full[14]), .A2(pipeline_csr_time_full[15]), .ZN(vscale_core_DW01_inc_6n136) );
  XOR2_X2 vscale_core_DW01_inc_6_U166 ( .A(vscale_core_DW01_inc_6n142), .B(vscale_core_DW01_inc_6n143), .Z(pipeline_csr_N726) );
  XNOR2_X2 vscale_core_DW01_inc_6_U171 ( .A(vscale_core_DW01_inc_6n148), .B(vscale_core_DW01_inc_6n147), .ZN(pipeline_csr_N725) );
  NAND2_X2 vscale_core_DW01_inc_6_U172 ( .A1(vscale_core_DW01_inc_6n152), .A2(vscale_core_DW01_inc_6n144), .ZN(vscale_core_DW01_inc_6n143) );
  NAND2_X2 vscale_core_DW01_inc_6_U174 ( .A1(pipeline_csr_time_full[12]), .A2(pipeline_csr_time_full[13]), .ZN(vscale_core_DW01_inc_6n145) );
  XNOR2_X2 vscale_core_DW01_inc_6_U177 ( .A(vscale_core_DW01_inc_6n152), .B(vscale_core_DW01_inc_6n151), .ZN(pipeline_csr_N724) );
  XNOR2_X2 vscale_core_DW01_inc_6_U182 ( .A(vscale_core_DW01_inc_6n158), .B(vscale_core_DW01_inc_6n157), .ZN(pipeline_csr_N723) );
  NAND2_X2 vscale_core_DW01_inc_6_U184 ( .A1(vscale_core_DW01_inc_6n170), .A2(vscale_core_DW01_inc_6n154), .ZN(vscale_core_DW01_inc_6n153) );
  NAND2_X2 vscale_core_DW01_inc_6_U186 ( .A1(pipeline_csr_time_full[10]), .A2(pipeline_csr_time_full[11]), .ZN(vscale_core_DW01_inc_6n155) );
  XOR2_X2 vscale_core_DW01_inc_6_U189 ( .A(vscale_core_DW01_inc_6n161), .B(vscale_core_DW01_inc_6n162), .Z(pipeline_csr_N722) );
  XOR2_X2 vscale_core_DW01_inc_6_U194 ( .A(vscale_core_DW01_inc_6n166), .B(vscale_core_DW01_inc_6n167), .Z(pipeline_csr_N721) );
  NAND2_X2 vscale_core_DW01_inc_6_U195 ( .A1(vscale_core_DW01_inc_6n170), .A2(vscale_core_DW01_inc_6n163), .ZN(vscale_core_DW01_inc_6n162) );
  NAND2_X2 vscale_core_DW01_inc_6_U197 ( .A1(pipeline_csr_time_full[8]), .A2(pipeline_csr_time_full[9]), .ZN(vscale_core_DW01_inc_6n164) );
  XNOR2_X2 vscale_core_DW01_inc_6_U200 ( .A(vscale_core_DW01_inc_6n170), .B(vscale_core_DW01_inc_6n169), .ZN(pipeline_csr_N720) );
  NAND2_X2 vscale_core_DW01_inc_6_U201 ( .A1(vscale_core_DW01_inc_6n170), .A2(pipeline_csr_time_full[8]), .ZN(vscale_core_DW01_inc_6n167) );
  XOR2_X2 vscale_core_DW01_inc_6_U204 ( .A(vscale_core_DW01_inc_6n175), .B(vscale_core_DW01_inc_6n176), .Z(pipeline_csr_N719) );
  NAND2_X2 vscale_core_DW01_inc_6_U206 ( .A1(vscale_core_DW01_inc_6n172), .A2(vscale_core_DW01_inc_6n188), .ZN(vscale_core_DW01_inc_6n171) );
  NAND2_X2 vscale_core_DW01_inc_6_U208 ( .A1(pipeline_csr_time_full[6]), .A2(pipeline_csr_time_full[7]), .ZN(vscale_core_DW01_inc_6n173) );
  XNOR2_X2 vscale_core_DW01_inc_6_U211 ( .A(vscale_core_DW01_inc_6n179), .B(vscale_core_DW01_inc_6n178), .ZN(pipeline_csr_N718) );
  NAND2_X2 vscale_core_DW01_inc_6_U212 ( .A1(vscale_core_DW01_inc_6n179), .A2(pipeline_csr_time_full[6]), .ZN(vscale_core_DW01_inc_6n176) );
  XNOR2_X2 vscale_core_DW01_inc_6_U215 ( .A(vscale_core_DW01_inc_6n183), .B(vscale_core_DW01_inc_6n182), .ZN(pipeline_csr_N717) );
  NAND2_X2 vscale_core_DW01_inc_6_U217 ( .A1(pipeline_csr_time_full[4]), .A2(pipeline_csr_time_full[5]), .ZN(vscale_core_DW01_inc_6n180) );
  XOR2_X2 vscale_core_DW01_inc_6_U220 ( .A(vscale_core_DW01_inc_6n186), .B(vscale_core_DW01_inc_6n187), .Z(pipeline_csr_N716) );
  XOR2_X2 vscale_core_DW01_inc_6_U225 ( .A(vscale_core_DW01_inc_6n191), .B(vscale_core_DW01_inc_6n192), .Z(pipeline_csr_N715) );
  NAND2_X2 vscale_core_DW01_inc_6_U228 ( .A1(pipeline_csr_time_full[2]), .A2(pipeline_csr_time_full[3]), .ZN(vscale_core_DW01_inc_6n189) );
  XNOR2_X2 vscale_core_DW01_inc_6_U231 ( .A(vscale_core_DW01_inc_6n195), .B(vscale_core_DW01_inc_6n194), .ZN(pipeline_csr_N714) );
  NAND2_X2 vscale_core_DW01_inc_6_U232 ( .A1(vscale_core_DW01_inc_6n195), .A2(pipeline_csr_time_full[2]), .ZN(vscale_core_DW01_inc_6n192) );
  XNOR2_X2 vscale_core_DW01_inc_6_U235 ( .A(vscale_core_DW01_inc_6n198), .B(pipeline_csr_time_full[0]), .ZN(pipeline_csr_N713) );
  NAND2_X2 vscale_core_DW01_inc_6_U237 ( .A1(pipeline_csr_time_full[1]), .A2(pipeline_csr_time_full[0]), .ZN(vscale_core_DW01_inc_6n196) );
  NOR2_X2 vscale_core_DW01_inc_6_U244 ( .A1(vscale_core_DW01_inc_6n99), .A2(vscale_core_DW01_inc_6n65), .ZN(vscale_core_DW01_inc_6n64) );
  NOR2_X2 vscale_core_DW01_inc_6_U245 ( .A1(vscale_core_DW01_inc_6n74), .A2(vscale_core_DW01_inc_6n67), .ZN(vscale_core_DW01_inc_6n66) );
  NOR2_X2 vscale_core_DW01_inc_6_U246 ( .A1(vscale_core_DW01_inc_6n37), .A2(vscale_core_DW01_inc_6n34), .ZN(vscale_core_DW01_inc_6n33) );
  NOR2_X2 vscale_core_DW01_inc_6_U247 ( .A1(vscale_core_DW01_inc_6n32), .A2(vscale_core_DW01_inc_6n29), .ZN(vscale_core_DW01_inc_6n28) );
  NOR2_X2 vscale_core_DW01_inc_6_U248 ( .A1(vscale_core_DW01_inc_6n132), .A2(vscale_core_DW01_inc_6n99), .ZN(vscale_core_DW01_inc_6n98) );
  NOR2_X2 vscale_core_DW01_inc_6_U249 ( .A1(vscale_core_DW01_inc_6n132), .A2(vscale_core_DW01_inc_6n116), .ZN(vscale_core_DW01_inc_6n115) );
  NOR2_X2 vscale_core_DW01_inc_6_U250 ( .A1(vscale_core_DW01_inc_6n97), .A2(vscale_core_DW01_inc_6n82), .ZN(vscale_core_DW01_inc_6n81) );
  NOR2_X2 vscale_core_DW01_inc_6_U251 ( .A1(vscale_core_DW01_inc_6n97), .A2(vscale_core_DW01_inc_6n91), .ZN(vscale_core_DW01_inc_6n90) );
  NOR2_X2 vscale_core_DW01_inc_6_U252 ( .A1(vscale_core_DW01_inc_6n80), .A2(vscale_core_DW01_inc_6n74), .ZN(vscale_core_DW01_inc_6n73) );
  NOR2_X2 vscale_core_DW01_inc_6_U253 ( .A1(vscale_core_DW01_inc_6n114), .A2(vscale_core_DW01_inc_6n108), .ZN(vscale_core_DW01_inc_6n107) );
  NOR2_X2 vscale_core_DW01_inc_6_U254 ( .A1(vscale_core_DW01_inc_6n132), .A2(vscale_core_DW01_inc_6n125), .ZN(vscale_core_DW01_inc_6n124) );
  NOR2_X2 vscale_core_DW01_inc_6_U255 ( .A1(vscale_core_DW01_inc_6n187), .A2(vscale_core_DW01_inc_6n180), .ZN(vscale_core_DW01_inc_6n179) );
  NOR2_X2 vscale_core_DW01_inc_6_U256 ( .A1(vscale_core_DW01_inc_6n132), .A2(vscale_core_DW01_inc_6n131), .ZN(vscale_core_DW01_inc_6n128) );
  NOR2_X2 vscale_core_DW01_inc_6_U257 ( .A1(vscale_core_DW01_inc_6n143), .A2(vscale_core_DW01_inc_6n142), .ZN(vscale_core_DW01_inc_6n139) );
  NOR2_X2 vscale_core_DW01_inc_6_U258 ( .A1(vscale_core_DW01_inc_6n153), .A2(vscale_core_DW01_inc_6n151), .ZN(vscale_core_DW01_inc_6n148) );
  NOR2_X2 vscale_core_DW01_inc_6_U259 ( .A1(vscale_core_DW01_inc_6n162), .A2(vscale_core_DW01_inc_6n161), .ZN(vscale_core_DW01_inc_6n158) );
  NOR2_X2 vscale_core_DW01_inc_6_U260 ( .A1(vscale_core_DW01_inc_6n45), .A2(vscale_core_DW01_inc_6n43), .ZN(vscale_core_DW01_inc_6n40) );
  NOR2_X2 vscale_core_DW01_inc_6_U261 ( .A1(vscale_core_DW01_inc_6n54), .A2(vscale_core_DW01_inc_6n53), .ZN(vscale_core_DW01_inc_6n50) );
  NOR2_X2 vscale_core_DW01_inc_6_U262 ( .A1(vscale_core_DW01_inc_6n187), .A2(vscale_core_DW01_inc_6n186), .ZN(vscale_core_DW01_inc_6n183) );
  NOR2_X2 vscale_core_DW01_inc_6_U263 ( .A1(vscale_core_DW01_inc_6n108), .A2(vscale_core_DW01_inc_6n101), .ZN(vscale_core_DW01_inc_6n100) );
  NOR2_X2 vscale_core_DW01_inc_6_U264 ( .A1(vscale_core_DW01_inc_6n180), .A2(vscale_core_DW01_inc_6n173), .ZN(vscale_core_DW01_inc_6n172) );
  NOR2_X2 vscale_core_DW01_inc_6_U265 ( .A1(vscale_core_DW01_inc_6n125), .A2(vscale_core_DW01_inc_6n118), .ZN(vscale_core_DW01_inc_6n117) );
  NOR2_X2 vscale_core_DW01_inc_6_U266 ( .A1(vscale_core_DW01_inc_6n91), .A2(vscale_core_DW01_inc_6n84), .ZN(vscale_core_DW01_inc_6n83) );
  NOR2_X2 vscale_core_DW01_inc_6_U267 ( .A1(vscale_core_DW01_inc_6n189), .A2(vscale_core_DW01_inc_6n196), .ZN(vscale_core_DW01_inc_6n188) );
  NOR2_X2 vscale_core_DW01_inc_6_U268 ( .A1(vscale_core_DW01_inc_6n134), .A2(vscale_core_DW01_inc_6n171), .ZN(vscale_core_DW01_inc_6n133) );
  NOR2_X2 vscale_core_DW01_inc_6_U269 ( .A1(vscale_core_DW01_inc_6n145), .A2(vscale_core_DW01_inc_6n136), .ZN(vscale_core_DW01_inc_6n135) );
  NOR2_X2 vscale_core_DW01_inc_6_U270 ( .A1(vscale_core_DW01_inc_6n164), .A2(vscale_core_DW01_inc_6n155), .ZN(vscale_core_DW01_inc_6n154) );
  NOR2_X2 vscale_core_DW01_inc_6_U271 ( .A1(vscale_core_DW01_inc_6n63), .A2(vscale_core_DW01_inc_6n24), .ZN(vscale_core_DW01_inc_6n23) );
  NOR2_X2 vscale_core_DW01_inc_6_U272 ( .A1(vscale_core_DW01_inc_6n56), .A2(vscale_core_DW01_inc_6n47), .ZN(vscale_core_DW01_inc_6n46) );
  INV_X4 vscale_core_DW01_inc_6_U273 ( .A(vscale_core_DW01_inc_6n98), .ZN(vscale_core_DW01_inc_6n97) );
  INV_X4 vscale_core_DW01_inc_6_U274 ( .A(pipeline_csr_time_full[24]), .ZN(vscale_core_DW01_inc_6n96) );
  INV_X4 vscale_core_DW01_inc_6_U275 ( .A(pipeline_csr_time_full[25]), .ZN(vscale_core_DW01_inc_6n93) );
  INV_X4 vscale_core_DW01_inc_6_U276 ( .A(pipeline_csr_time_full[26]), .ZN(vscale_core_DW01_inc_6n89) );
  INV_X4 vscale_core_DW01_inc_6_U277 ( .A(pipeline_csr_time_full[27]), .ZN(vscale_core_DW01_inc_6n86) );
  INV_X4 vscale_core_DW01_inc_6_U278 ( .A(vscale_core_DW01_inc_6n83), .ZN(vscale_core_DW01_inc_6n82) );
  INV_X4 vscale_core_DW01_inc_6_U279 ( .A(vscale_core_DW01_inc_6n81), .ZN(vscale_core_DW01_inc_6n80) );
  INV_X4 vscale_core_DW01_inc_6_U280 ( .A(pipeline_csr_time_full[28]), .ZN(vscale_core_DW01_inc_6n79) );
  INV_X4 vscale_core_DW01_inc_6_U281 ( .A(pipeline_csr_time_full[29]), .ZN(vscale_core_DW01_inc_6n76) );
  INV_X4 vscale_core_DW01_inc_6_U282 ( .A(pipeline_csr_time_full[30]), .ZN(vscale_core_DW01_inc_6n72) );
  INV_X4 vscale_core_DW01_inc_6_U283 ( .A(pipeline_csr_time_full[31]), .ZN(vscale_core_DW01_inc_6n69) );
  INV_X4 vscale_core_DW01_inc_6_U284 ( .A(vscale_core_DW01_inc_6n63), .ZN(vscale_core_DW01_inc_6n62) );
  INV_X4 vscale_core_DW01_inc_6_U285 ( .A(pipeline_csr_time_full[32]), .ZN(vscale_core_DW01_inc_6n61) );
  INV_X4 vscale_core_DW01_inc_6_U286 ( .A(pipeline_csr_time_full[33]), .ZN(vscale_core_DW01_inc_6n58) );
  INV_X4 vscale_core_DW01_inc_6_U287 ( .A(vscale_core_DW01_inc_6n56), .ZN(vscale_core_DW01_inc_6n55) );
  INV_X4 vscale_core_DW01_inc_6_U288 ( .A(pipeline_csr_time_full[34]), .ZN(vscale_core_DW01_inc_6n53) );
  INV_X4 vscale_core_DW01_inc_6_U289 ( .A(pipeline_csr_time_full[35]), .ZN(vscale_core_DW01_inc_6n49) );
  INV_X4 vscale_core_DW01_inc_6_U290 ( .A(vscale_core_DW01_inc_6n45), .ZN(vscale_core_DW01_inc_6n44) );
  INV_X4 vscale_core_DW01_inc_6_U291 ( .A(pipeline_csr_time_full[36]), .ZN(vscale_core_DW01_inc_6n43) );
  INV_X4 vscale_core_DW01_inc_6_U292 ( .A(pipeline_csr_time_full[37]), .ZN(vscale_core_DW01_inc_6n39) );
  INV_X4 vscale_core_DW01_inc_6_U293 ( .A(vscale_core_DW01_inc_6n37), .ZN(vscale_core_DW01_inc_6n36) );
  INV_X4 vscale_core_DW01_inc_6_U294 ( .A(pipeline_csr_time_full[38]), .ZN(vscale_core_DW01_inc_6n34) );
  INV_X4 vscale_core_DW01_inc_6_U295 ( .A(vscale_core_DW01_inc_6n32), .ZN(vscale_core_DW01_inc_6n31) );
  INV_X4 vscale_core_DW01_inc_6_U296 ( .A(pipeline_csr_time_full[39]), .ZN(vscale_core_DW01_inc_6n29) );
  INV_X4 vscale_core_DW01_inc_6_U297 ( .A(pipeline_csr_time_full[40]), .ZN(vscale_core_DW01_inc_6n26) );
  INV_X4 vscale_core_DW01_inc_6_U298 ( .A(pipeline_csr_time_full[1]), .ZN(vscale_core_DW01_inc_6n198) );
  INV_X4 vscale_core_DW01_inc_6_U299 ( .A(vscale_core_DW01_inc_6n196), .ZN(vscale_core_DW01_inc_6n195) );
  INV_X4 vscale_core_DW01_inc_6_U300 ( .A(pipeline_csr_time_full[2]), .ZN(vscale_core_DW01_inc_6n194) );
  INV_X4 vscale_core_DW01_inc_6_U301 ( .A(pipeline_csr_time_full[3]), .ZN(vscale_core_DW01_inc_6n191) );
  INV_X4 vscale_core_DW01_inc_6_U302 ( .A(vscale_core_DW01_inc_6n188), .ZN(vscale_core_DW01_inc_6n187) );
  INV_X4 vscale_core_DW01_inc_6_U303 ( .A(pipeline_csr_time_full[4]), .ZN(vscale_core_DW01_inc_6n186) );
  INV_X4 vscale_core_DW01_inc_6_U304 ( .A(pipeline_csr_time_full[5]), .ZN(vscale_core_DW01_inc_6n182) );
  INV_X4 vscale_core_DW01_inc_6_U305 ( .A(pipeline_csr_time_full[6]), .ZN(vscale_core_DW01_inc_6n178) );
  INV_X4 vscale_core_DW01_inc_6_U306 ( .A(pipeline_csr_time_full[7]), .ZN(vscale_core_DW01_inc_6n175) );
  INV_X4 vscale_core_DW01_inc_6_U307 ( .A(vscale_core_DW01_inc_6n171), .ZN(vscale_core_DW01_inc_6n170) );
  INV_X4 vscale_core_DW01_inc_6_U308 ( .A(pipeline_csr_time_full[8]), .ZN(vscale_core_DW01_inc_6n169) );
  INV_X4 vscale_core_DW01_inc_6_U309 ( .A(pipeline_csr_time_full[9]), .ZN(vscale_core_DW01_inc_6n166) );
  INV_X4 vscale_core_DW01_inc_6_U310 ( .A(vscale_core_DW01_inc_6n164), .ZN(vscale_core_DW01_inc_6n163) );
  INV_X4 vscale_core_DW01_inc_6_U311 ( .A(pipeline_csr_time_full[10]), .ZN(vscale_core_DW01_inc_6n161) );
  INV_X4 vscale_core_DW01_inc_6_U312 ( .A(pipeline_csr_time_full[11]), .ZN(vscale_core_DW01_inc_6n157) );
  INV_X4 vscale_core_DW01_inc_6_U313 ( .A(vscale_core_DW01_inc_6n153), .ZN(vscale_core_DW01_inc_6n152) );
  INV_X4 vscale_core_DW01_inc_6_U314 ( .A(pipeline_csr_time_full[12]), .ZN(vscale_core_DW01_inc_6n151) );
  INV_X4 vscale_core_DW01_inc_6_U315 ( .A(pipeline_csr_time_full[13]), .ZN(vscale_core_DW01_inc_6n147) );
  INV_X4 vscale_core_DW01_inc_6_U316 ( .A(vscale_core_DW01_inc_6n145), .ZN(vscale_core_DW01_inc_6n144) );
  INV_X4 vscale_core_DW01_inc_6_U317 ( .A(pipeline_csr_time_full[14]), .ZN(vscale_core_DW01_inc_6n142) );
  INV_X4 vscale_core_DW01_inc_6_U318 ( .A(pipeline_csr_time_full[15]), .ZN(vscale_core_DW01_inc_6n138) );
  INV_X4 vscale_core_DW01_inc_6_U319 ( .A(vscale_core_DW01_inc_6n133), .ZN(vscale_core_DW01_inc_6n132) );
  INV_X4 vscale_core_DW01_inc_6_U320 ( .A(pipeline_csr_time_full[16]), .ZN(vscale_core_DW01_inc_6n131) );
  INV_X4 vscale_core_DW01_inc_6_U321 ( .A(pipeline_csr_time_full[17]), .ZN(vscale_core_DW01_inc_6n127) );
  INV_X4 vscale_core_DW01_inc_6_U322 ( .A(pipeline_csr_time_full[18]), .ZN(vscale_core_DW01_inc_6n123) );
  INV_X4 vscale_core_DW01_inc_6_U323 ( .A(pipeline_csr_time_full[19]), .ZN(vscale_core_DW01_inc_6n120) );
  INV_X4 vscale_core_DW01_inc_6_U324 ( .A(vscale_core_DW01_inc_6n117), .ZN(vscale_core_DW01_inc_6n116) );
  INV_X4 vscale_core_DW01_inc_6_U325 ( .A(vscale_core_DW01_inc_6n115), .ZN(vscale_core_DW01_inc_6n114) );
  INV_X4 vscale_core_DW01_inc_6_U326 ( .A(pipeline_csr_time_full[20]), .ZN(vscale_core_DW01_inc_6n113) );
  INV_X4 vscale_core_DW01_inc_6_U327 ( .A(pipeline_csr_time_full[21]), .ZN(vscale_core_DW01_inc_6n110) );
  INV_X4 vscale_core_DW01_inc_6_U328 ( .A(pipeline_csr_time_full[22]), .ZN(vscale_core_DW01_inc_6n106) );
  INV_X4 vscale_core_DW01_inc_6_U329 ( .A(pipeline_csr_time_full[23]), .ZN(vscale_core_DW01_inc_6n103) );
  INV_X4 vscale_core_DW01_inc_6_U330 ( .A(pipeline_csr_time_full[0]), .ZN(pipeline_csr_N712) );
;
  vscale_core_DW01_inc_7 pipeline_csr_add_311 

  XOR2_X2 vscale_core_DW01_inc_7_U1 ( .A(pipeline_csr_cycle_full[63]), .B(vscale_core_DW01_inc_7n1), .Z(pipeline_csr_N711) );
  HA_X1 vscale_core_DW01_inc_7_U2 ( .A(pipeline_csr_cycle_full[62]), .B(vscale_core_DW01_inc_7n2), .CO(vscale_core_DW01_inc_7n1), .S(pipeline_csr_N710) );
  HA_X1 vscale_core_DW01_inc_7_U3 ( .A(pipeline_csr_cycle_full[61]), .B(vscale_core_DW01_inc_7n3), .CO(vscale_core_DW01_inc_7n2), .S(pipeline_csr_N709) );
  HA_X1 vscale_core_DW01_inc_7_U4 ( .A(pipeline_csr_cycle_full[60]), .B(vscale_core_DW01_inc_7n4), .CO(vscale_core_DW01_inc_7n3), .S(pipeline_csr_N708) );
  HA_X1 vscale_core_DW01_inc_7_U5 ( .A(pipeline_csr_cycle_full[59]), .B(vscale_core_DW01_inc_7n5), .CO(vscale_core_DW01_inc_7n4), .S(pipeline_csr_N707) );
  HA_X1 vscale_core_DW01_inc_7_U6 ( .A(pipeline_csr_cycle_full[58]), .B(vscale_core_DW01_inc_7n6), .CO(vscale_core_DW01_inc_7n5), .S(pipeline_csr_N706) );
  HA_X1 vscale_core_DW01_inc_7_U7 ( .A(pipeline_csr_cycle_full[57]), .B(vscale_core_DW01_inc_7n7), .CO(vscale_core_DW01_inc_7n6), .S(pipeline_csr_N705) );
  HA_X1 vscale_core_DW01_inc_7_U8 ( .A(pipeline_csr_cycle_full[56]), .B(vscale_core_DW01_inc_7n8), .CO(vscale_core_DW01_inc_7n7), .S(pipeline_csr_N704) );
  HA_X1 vscale_core_DW01_inc_7_U9 ( .A(pipeline_csr_cycle_full[55]), .B(vscale_core_DW01_inc_7n9), .CO(vscale_core_DW01_inc_7n8), .S(pipeline_csr_N703) );
  HA_X1 vscale_core_DW01_inc_7_U10 ( .A(pipeline_csr_cycle_full[54]), .B(vscale_core_DW01_inc_7n10), .CO(vscale_core_DW01_inc_7n9), .S(pipeline_csr_N702) );
  HA_X1 vscale_core_DW01_inc_7_U11 ( .A(pipeline_csr_cycle_full[53]), .B(vscale_core_DW01_inc_7n11), .CO(vscale_core_DW01_inc_7n10), .S(pipeline_csr_N701) );
  HA_X1 vscale_core_DW01_inc_7_U12 ( .A(pipeline_csr_cycle_full[52]), .B(vscale_core_DW01_inc_7n12), .CO(vscale_core_DW01_inc_7n11), .S(pipeline_csr_N700) );
  HA_X1 vscale_core_DW01_inc_7_U13 ( .A(pipeline_csr_cycle_full[51]), .B(vscale_core_DW01_inc_7n13), .CO(vscale_core_DW01_inc_7n12), .S(pipeline_csr_N699) );
  HA_X1 vscale_core_DW01_inc_7_U14 ( .A(pipeline_csr_cycle_full[50]), .B(vscale_core_DW01_inc_7n14), .CO(vscale_core_DW01_inc_7n13), .S(pipeline_csr_N698) );
  HA_X1 vscale_core_DW01_inc_7_U15 ( .A(pipeline_csr_cycle_full[49]), .B(vscale_core_DW01_inc_7n15), .CO(vscale_core_DW01_inc_7n14), .S(pipeline_csr_N697) );
  HA_X1 vscale_core_DW01_inc_7_U16 ( .A(pipeline_csr_cycle_full[48]), .B(vscale_core_DW01_inc_7n16), .CO(vscale_core_DW01_inc_7n15), .S(pipeline_csr_N696) );
  HA_X1 vscale_core_DW01_inc_7_U17 ( .A(pipeline_csr_cycle_full[47]), .B(vscale_core_DW01_inc_7n17), .CO(vscale_core_DW01_inc_7n16), .S(pipeline_csr_N695) );
  HA_X1 vscale_core_DW01_inc_7_U18 ( .A(pipeline_csr_cycle_full[46]), .B(vscale_core_DW01_inc_7n18), .CO(vscale_core_DW01_inc_7n17), .S(pipeline_csr_N694) );
  HA_X1 vscale_core_DW01_inc_7_U19 ( .A(pipeline_csr_cycle_full[45]), .B(vscale_core_DW01_inc_7n19), .CO(vscale_core_DW01_inc_7n18), .S(pipeline_csr_N693) );
  HA_X1 vscale_core_DW01_inc_7_U20 ( .A(pipeline_csr_cycle_full[44]), .B(vscale_core_DW01_inc_7n20), .CO(vscale_core_DW01_inc_7n19), .S(pipeline_csr_N692) );
  HA_X1 vscale_core_DW01_inc_7_U21 ( .A(pipeline_csr_cycle_full[43]), .B(vscale_core_DW01_inc_7n21), .CO(vscale_core_DW01_inc_7n20), .S(pipeline_csr_N691) );
  HA_X1 vscale_core_DW01_inc_7_U22 ( .A(pipeline_csr_cycle_full[42]), .B(vscale_core_DW01_inc_7n22), .CO(vscale_core_DW01_inc_7n21), .S(pipeline_csr_N690) );
  HA_X1 vscale_core_DW01_inc_7_U23 ( .A(pipeline_csr_cycle_full[41]), .B(vscale_core_DW01_inc_7n23), .CO(vscale_core_DW01_inc_7n22), .S(pipeline_csr_N689) );
  XOR2_X2 vscale_core_DW01_inc_7_U24 ( .A(vscale_core_DW01_inc_7n26), .B(vscale_core_DW01_inc_7n27), .Z(pipeline_csr_N688) );
  NAND2_X2 vscale_core_DW01_inc_7_U26 ( .A1(vscale_core_DW01_inc_7n28), .A2(pipeline_csr_cycle_full[40]), .ZN(vscale_core_DW01_inc_7n24) );
  XOR2_X2 vscale_core_DW01_inc_7_U29 ( .A(vscale_core_DW01_inc_7n29), .B(vscale_core_DW01_inc_7n30), .Z(pipeline_csr_N687) );
  NAND2_X2 vscale_core_DW01_inc_7_U30 ( .A1(vscale_core_DW01_inc_7n62), .A2(vscale_core_DW01_inc_7n28), .ZN(vscale_core_DW01_inc_7n27) );
  XOR2_X2 vscale_core_DW01_inc_7_U33 ( .A(vscale_core_DW01_inc_7n34), .B(vscale_core_DW01_inc_7n35), .Z(pipeline_csr_N686) );
  NAND2_X2 vscale_core_DW01_inc_7_U34 ( .A1(vscale_core_DW01_inc_7n62), .A2(vscale_core_DW01_inc_7n31), .ZN(vscale_core_DW01_inc_7n30) );
  NAND2_X2 vscale_core_DW01_inc_7_U36 ( .A1(vscale_core_DW01_inc_7n46), .A2(vscale_core_DW01_inc_7n33), .ZN(vscale_core_DW01_inc_7n32) );
  XNOR2_X2 vscale_core_DW01_inc_7_U39 ( .A(vscale_core_DW01_inc_7n40), .B(vscale_core_DW01_inc_7n39), .ZN(pipeline_csr_N685) );
  NAND2_X2 vscale_core_DW01_inc_7_U40 ( .A1(vscale_core_DW01_inc_7n44), .A2(vscale_core_DW01_inc_7n36), .ZN(vscale_core_DW01_inc_7n35) );
  NAND2_X2 vscale_core_DW01_inc_7_U42 ( .A1(pipeline_csr_cycle_full[36]), .A2(pipeline_csr_cycle_full[37]), .ZN(vscale_core_DW01_inc_7n37) );
  XNOR2_X2 vscale_core_DW01_inc_7_U45 ( .A(vscale_core_DW01_inc_7n44), .B(vscale_core_DW01_inc_7n43), .ZN(pipeline_csr_N684) );
  XNOR2_X2 vscale_core_DW01_inc_7_U50 ( .A(vscale_core_DW01_inc_7n50), .B(vscale_core_DW01_inc_7n49), .ZN(pipeline_csr_N683) );
  NAND2_X2 vscale_core_DW01_inc_7_U52 ( .A1(vscale_core_DW01_inc_7n62), .A2(vscale_core_DW01_inc_7n46), .ZN(vscale_core_DW01_inc_7n45) );
  NAND2_X2 vscale_core_DW01_inc_7_U54 ( .A1(pipeline_csr_cycle_full[34]), .A2(pipeline_csr_cycle_full[35]), .ZN(vscale_core_DW01_inc_7n47) );
  XOR2_X2 vscale_core_DW01_inc_7_U57 ( .A(vscale_core_DW01_inc_7n53), .B(vscale_core_DW01_inc_7n54), .Z(pipeline_csr_N682) );
  XOR2_X2 vscale_core_DW01_inc_7_U62 ( .A(vscale_core_DW01_inc_7n58), .B(vscale_core_DW01_inc_7n59), .Z(pipeline_csr_N681) );
  NAND2_X2 vscale_core_DW01_inc_7_U63 ( .A1(vscale_core_DW01_inc_7n62), .A2(vscale_core_DW01_inc_7n55), .ZN(vscale_core_DW01_inc_7n54) );
  NAND2_X2 vscale_core_DW01_inc_7_U65 ( .A1(pipeline_csr_cycle_full[32]), .A2(pipeline_csr_cycle_full[33]), .ZN(vscale_core_DW01_inc_7n56) );
  XNOR2_X2 vscale_core_DW01_inc_7_U68 ( .A(vscale_core_DW01_inc_7n62), .B(vscale_core_DW01_inc_7n61), .ZN(pipeline_csr_N680) );
  NAND2_X2 vscale_core_DW01_inc_7_U69 ( .A1(vscale_core_DW01_inc_7n62), .A2(pipeline_csr_cycle_full[32]), .ZN(vscale_core_DW01_inc_7n59) );
  XOR2_X2 vscale_core_DW01_inc_7_U72 ( .A(vscale_core_DW01_inc_7n69), .B(vscale_core_DW01_inc_7n70), .Z(pipeline_csr_N679) );
  NAND2_X2 vscale_core_DW01_inc_7_U74 ( .A1(vscale_core_DW01_inc_7n64), .A2(vscale_core_DW01_inc_7n133), .ZN(vscale_core_DW01_inc_7n63) );
  NAND2_X2 vscale_core_DW01_inc_7_U76 ( .A1(vscale_core_DW01_inc_7n83), .A2(vscale_core_DW01_inc_7n66), .ZN(vscale_core_DW01_inc_7n65) );
  NAND2_X2 vscale_core_DW01_inc_7_U78 ( .A1(pipeline_csr_cycle_full[30]), .A2(pipeline_csr_cycle_full[31]), .ZN(vscale_core_DW01_inc_7n67) );
  XNOR2_X2 vscale_core_DW01_inc_7_U81 ( .A(vscale_core_DW01_inc_7n73), .B(vscale_core_DW01_inc_7n72), .ZN(pipeline_csr_N678) );
  NAND2_X2 vscale_core_DW01_inc_7_U82 ( .A1(vscale_core_DW01_inc_7n73), .A2(pipeline_csr_cycle_full[30]), .ZN(vscale_core_DW01_inc_7n70) );
  XOR2_X2 vscale_core_DW01_inc_7_U85 ( .A(vscale_core_DW01_inc_7n76), .B(vscale_core_DW01_inc_7n77), .Z(pipeline_csr_N677) );
  NAND2_X2 vscale_core_DW01_inc_7_U87 ( .A1(pipeline_csr_cycle_full[28]), .A2(pipeline_csr_cycle_full[29]), .ZN(vscale_core_DW01_inc_7n74) );
  XOR2_X2 vscale_core_DW01_inc_7_U90 ( .A(vscale_core_DW01_inc_7n79), .B(vscale_core_DW01_inc_7n80), .Z(pipeline_csr_N676) );
  NAND2_X2 vscale_core_DW01_inc_7_U91 ( .A1(vscale_core_DW01_inc_7n81), .A2(pipeline_csr_cycle_full[28]), .ZN(vscale_core_DW01_inc_7n77) );
  XOR2_X2 vscale_core_DW01_inc_7_U94 ( .A(vscale_core_DW01_inc_7n86), .B(vscale_core_DW01_inc_7n87), .Z(pipeline_csr_N675) );
  NAND2_X2 vscale_core_DW01_inc_7_U99 ( .A1(pipeline_csr_cycle_full[26]), .A2(pipeline_csr_cycle_full[27]), .ZN(vscale_core_DW01_inc_7n84) );
  XNOR2_X2 vscale_core_DW01_inc_7_U102 ( .A(vscale_core_DW01_inc_7n90), .B(vscale_core_DW01_inc_7n89), .ZN(pipeline_csr_N674) );
  NAND2_X2 vscale_core_DW01_inc_7_U103 ( .A1(vscale_core_DW01_inc_7n90), .A2(pipeline_csr_cycle_full[26]), .ZN(vscale_core_DW01_inc_7n87) );
  XOR2_X2 vscale_core_DW01_inc_7_U106 ( .A(vscale_core_DW01_inc_7n93), .B(vscale_core_DW01_inc_7n94), .Z(pipeline_csr_N673) );
  NAND2_X2 vscale_core_DW01_inc_7_U108 ( .A1(pipeline_csr_cycle_full[24]), .A2(pipeline_csr_cycle_full[25]), .ZN(vscale_core_DW01_inc_7n91) );
  XOR2_X2 vscale_core_DW01_inc_7_U111 ( .A(vscale_core_DW01_inc_7n96), .B(vscale_core_DW01_inc_7n97), .Z(pipeline_csr_N672) );
  NAND2_X2 vscale_core_DW01_inc_7_U112 ( .A1(vscale_core_DW01_inc_7n98), .A2(pipeline_csr_cycle_full[24]), .ZN(vscale_core_DW01_inc_7n94) );
  XOR2_X2 vscale_core_DW01_inc_7_U115 ( .A(vscale_core_DW01_inc_7n103), .B(vscale_core_DW01_inc_7n104), .Z(pipeline_csr_N671) );
  NAND2_X2 vscale_core_DW01_inc_7_U118 ( .A1(vscale_core_DW01_inc_7n117), .A2(vscale_core_DW01_inc_7n100), .ZN(vscale_core_DW01_inc_7n99) );
  NAND2_X2 vscale_core_DW01_inc_7_U120 ( .A1(pipeline_csr_cycle_full[22]), .A2(pipeline_csr_cycle_full[23]), .ZN(vscale_core_DW01_inc_7n101) );
  XNOR2_X2 vscale_core_DW01_inc_7_U123 ( .A(vscale_core_DW01_inc_7n107), .B(vscale_core_DW01_inc_7n106), .ZN(pipeline_csr_N670) );
  NAND2_X2 vscale_core_DW01_inc_7_U124 ( .A1(vscale_core_DW01_inc_7n107), .A2(pipeline_csr_cycle_full[22]), .ZN(vscale_core_DW01_inc_7n104) );
  XOR2_X2 vscale_core_DW01_inc_7_U127 ( .A(vscale_core_DW01_inc_7n110), .B(vscale_core_DW01_inc_7n111), .Z(pipeline_csr_N669) );
  NAND2_X2 vscale_core_DW01_inc_7_U129 ( .A1(pipeline_csr_cycle_full[20]), .A2(pipeline_csr_cycle_full[21]), .ZN(vscale_core_DW01_inc_7n108) );
  XOR2_X2 vscale_core_DW01_inc_7_U132 ( .A(vscale_core_DW01_inc_7n113), .B(vscale_core_DW01_inc_7n114), .Z(pipeline_csr_N668) );
  NAND2_X2 vscale_core_DW01_inc_7_U133 ( .A1(vscale_core_DW01_inc_7n115), .A2(pipeline_csr_cycle_full[20]), .ZN(vscale_core_DW01_inc_7n111) );
  XOR2_X2 vscale_core_DW01_inc_7_U136 ( .A(vscale_core_DW01_inc_7n120), .B(vscale_core_DW01_inc_7n121), .Z(pipeline_csr_N667) );
  NAND2_X2 vscale_core_DW01_inc_7_U141 ( .A1(pipeline_csr_cycle_full[18]), .A2(pipeline_csr_cycle_full[19]), .ZN(vscale_core_DW01_inc_7n118) );
  XNOR2_X2 vscale_core_DW01_inc_7_U144 ( .A(vscale_core_DW01_inc_7n124), .B(vscale_core_DW01_inc_7n123), .ZN(pipeline_csr_N666) );
  NAND2_X2 vscale_core_DW01_inc_7_U145 ( .A1(vscale_core_DW01_inc_7n124), .A2(pipeline_csr_cycle_full[18]), .ZN(vscale_core_DW01_inc_7n121) );
  XNOR2_X2 vscale_core_DW01_inc_7_U148 ( .A(vscale_core_DW01_inc_7n128), .B(vscale_core_DW01_inc_7n127), .ZN(pipeline_csr_N665) );
  NAND2_X2 vscale_core_DW01_inc_7_U150 ( .A1(pipeline_csr_cycle_full[16]), .A2(pipeline_csr_cycle_full[17]), .ZN(vscale_core_DW01_inc_7n125) );
  XOR2_X2 vscale_core_DW01_inc_7_U153 ( .A(vscale_core_DW01_inc_7n131), .B(vscale_core_DW01_inc_7n132), .Z(pipeline_csr_N664) );
  XNOR2_X2 vscale_core_DW01_inc_7_U158 ( .A(vscale_core_DW01_inc_7n139), .B(vscale_core_DW01_inc_7n138), .ZN(pipeline_csr_N663) );
  NAND2_X2 vscale_core_DW01_inc_7_U161 ( .A1(vscale_core_DW01_inc_7n154), .A2(vscale_core_DW01_inc_7n135), .ZN(vscale_core_DW01_inc_7n134) );
  NAND2_X2 vscale_core_DW01_inc_7_U163 ( .A1(pipeline_csr_cycle_full[14]), .A2(pipeline_csr_cycle_full[15]), .ZN(vscale_core_DW01_inc_7n136) );
  XOR2_X2 vscale_core_DW01_inc_7_U166 ( .A(vscale_core_DW01_inc_7n142), .B(vscale_core_DW01_inc_7n143), .Z(pipeline_csr_N662) );
  XNOR2_X2 vscale_core_DW01_inc_7_U171 ( .A(vscale_core_DW01_inc_7n148), .B(vscale_core_DW01_inc_7n147), .ZN(pipeline_csr_N661) );
  NAND2_X2 vscale_core_DW01_inc_7_U172 ( .A1(vscale_core_DW01_inc_7n152), .A2(vscale_core_DW01_inc_7n144), .ZN(vscale_core_DW01_inc_7n143) );
  NAND2_X2 vscale_core_DW01_inc_7_U174 ( .A1(pipeline_csr_cycle_full[12]), .A2(pipeline_csr_cycle_full[13]), .ZN(vscale_core_DW01_inc_7n145) );
  XNOR2_X2 vscale_core_DW01_inc_7_U177 ( .A(vscale_core_DW01_inc_7n152), .B(vscale_core_DW01_inc_7n151), .ZN(pipeline_csr_N660) );
  XNOR2_X2 vscale_core_DW01_inc_7_U182 ( .A(vscale_core_DW01_inc_7n158), .B(vscale_core_DW01_inc_7n157), .ZN(pipeline_csr_N659) );
  NAND2_X2 vscale_core_DW01_inc_7_U184 ( .A1(vscale_core_DW01_inc_7n170), .A2(vscale_core_DW01_inc_7n154), .ZN(vscale_core_DW01_inc_7n153) );
  NAND2_X2 vscale_core_DW01_inc_7_U186 ( .A1(pipeline_csr_cycle_full[10]), .A2(pipeline_csr_cycle_full[11]), .ZN(vscale_core_DW01_inc_7n155) );
  XOR2_X2 vscale_core_DW01_inc_7_U189 ( .A(vscale_core_DW01_inc_7n161), .B(vscale_core_DW01_inc_7n162), .Z(pipeline_csr_N658) );
  XOR2_X2 vscale_core_DW01_inc_7_U194 ( .A(vscale_core_DW01_inc_7n166), .B(vscale_core_DW01_inc_7n167), .Z(pipeline_csr_N657) );
  NAND2_X2 vscale_core_DW01_inc_7_U195 ( .A1(vscale_core_DW01_inc_7n170), .A2(vscale_core_DW01_inc_7n163), .ZN(vscale_core_DW01_inc_7n162) );
  NAND2_X2 vscale_core_DW01_inc_7_U197 ( .A1(pipeline_csr_cycle_full[8]), .A2(pipeline_csr_cycle_full[9]), .ZN(vscale_core_DW01_inc_7n164) );
  XNOR2_X2 vscale_core_DW01_inc_7_U200 ( .A(vscale_core_DW01_inc_7n170), .B(vscale_core_DW01_inc_7n169), .ZN(pipeline_csr_N656) );
  NAND2_X2 vscale_core_DW01_inc_7_U201 ( .A1(vscale_core_DW01_inc_7n170), .A2(pipeline_csr_cycle_full[8]), .ZN(vscale_core_DW01_inc_7n167) );
  XOR2_X2 vscale_core_DW01_inc_7_U204 ( .A(vscale_core_DW01_inc_7n175), .B(vscale_core_DW01_inc_7n176), .Z(pipeline_csr_N655) );
  NAND2_X2 vscale_core_DW01_inc_7_U206 ( .A1(vscale_core_DW01_inc_7n172), .A2(vscale_core_DW01_inc_7n188), .ZN(vscale_core_DW01_inc_7n171) );
  NAND2_X2 vscale_core_DW01_inc_7_U208 ( .A1(pipeline_csr_cycle_full[6]), .A2(pipeline_csr_cycle_full[7]), .ZN(vscale_core_DW01_inc_7n173) );
  XNOR2_X2 vscale_core_DW01_inc_7_U211 ( .A(vscale_core_DW01_inc_7n179), .B(vscale_core_DW01_inc_7n178), .ZN(pipeline_csr_N654) );
  NAND2_X2 vscale_core_DW01_inc_7_U212 ( .A1(vscale_core_DW01_inc_7n179), .A2(pipeline_csr_cycle_full[6]), .ZN(vscale_core_DW01_inc_7n176) );
  XNOR2_X2 vscale_core_DW01_inc_7_U215 ( .A(vscale_core_DW01_inc_7n183), .B(vscale_core_DW01_inc_7n182), .ZN(pipeline_csr_N653) );
  NAND2_X2 vscale_core_DW01_inc_7_U217 ( .A1(pipeline_csr_cycle_full[4]), .A2(pipeline_csr_cycle_full[5]), .ZN(vscale_core_DW01_inc_7n180) );
  XOR2_X2 vscale_core_DW01_inc_7_U220 ( .A(vscale_core_DW01_inc_7n186), .B(vscale_core_DW01_inc_7n187), .Z(pipeline_csr_N652) );
  XOR2_X2 vscale_core_DW01_inc_7_U225 ( .A(vscale_core_DW01_inc_7n191), .B(vscale_core_DW01_inc_7n192), .Z(pipeline_csr_N651) );
  NAND2_X2 vscale_core_DW01_inc_7_U228 ( .A1(pipeline_csr_cycle_full[2]), .A2(pipeline_csr_cycle_full[3]), .ZN(vscale_core_DW01_inc_7n189) );
  XNOR2_X2 vscale_core_DW01_inc_7_U231 ( .A(vscale_core_DW01_inc_7n195), .B(vscale_core_DW01_inc_7n194), .ZN(pipeline_csr_N650) );
  NAND2_X2 vscale_core_DW01_inc_7_U232 ( .A1(vscale_core_DW01_inc_7n195), .A2(pipeline_csr_cycle_full[2]), .ZN(vscale_core_DW01_inc_7n192) );
  XNOR2_X2 vscale_core_DW01_inc_7_U235 ( .A(vscale_core_DW01_inc_7n198), .B(pipeline_csr_cycle_full[0]), .ZN(pipeline_csr_N649) );
  NAND2_X2 vscale_core_DW01_inc_7_U237 ( .A1(pipeline_csr_cycle_full[1]), .A2(pipeline_csr_cycle_full[0]), .ZN(vscale_core_DW01_inc_7n196) );
  NOR2_X2 vscale_core_DW01_inc_7_U244 ( .A1(vscale_core_DW01_inc_7n99), .A2(vscale_core_DW01_inc_7n65), .ZN(vscale_core_DW01_inc_7n64) );
  NOR2_X2 vscale_core_DW01_inc_7_U245 ( .A1(vscale_core_DW01_inc_7n74), .A2(vscale_core_DW01_inc_7n67), .ZN(vscale_core_DW01_inc_7n66) );
  NOR2_X2 vscale_core_DW01_inc_7_U246 ( .A1(vscale_core_DW01_inc_7n37), .A2(vscale_core_DW01_inc_7n34), .ZN(vscale_core_DW01_inc_7n33) );
  NOR2_X2 vscale_core_DW01_inc_7_U247 ( .A1(vscale_core_DW01_inc_7n32), .A2(vscale_core_DW01_inc_7n29), .ZN(vscale_core_DW01_inc_7n28) );
  NOR2_X2 vscale_core_DW01_inc_7_U248 ( .A1(vscale_core_DW01_inc_7n132), .A2(vscale_core_DW01_inc_7n99), .ZN(vscale_core_DW01_inc_7n98) );
  NOR2_X2 vscale_core_DW01_inc_7_U249 ( .A1(vscale_core_DW01_inc_7n132), .A2(vscale_core_DW01_inc_7n116), .ZN(vscale_core_DW01_inc_7n115) );
  NOR2_X2 vscale_core_DW01_inc_7_U250 ( .A1(vscale_core_DW01_inc_7n97), .A2(vscale_core_DW01_inc_7n82), .ZN(vscale_core_DW01_inc_7n81) );
  NOR2_X2 vscale_core_DW01_inc_7_U251 ( .A1(vscale_core_DW01_inc_7n80), .A2(vscale_core_DW01_inc_7n74), .ZN(vscale_core_DW01_inc_7n73) );
  NOR2_X2 vscale_core_DW01_inc_7_U252 ( .A1(vscale_core_DW01_inc_7n114), .A2(vscale_core_DW01_inc_7n108), .ZN(vscale_core_DW01_inc_7n107) );
  NOR2_X2 vscale_core_DW01_inc_7_U253 ( .A1(vscale_core_DW01_inc_7n97), .A2(vscale_core_DW01_inc_7n91), .ZN(vscale_core_DW01_inc_7n90) );
  NOR2_X2 vscale_core_DW01_inc_7_U254 ( .A1(vscale_core_DW01_inc_7n132), .A2(vscale_core_DW01_inc_7n125), .ZN(vscale_core_DW01_inc_7n124) );
  NOR2_X2 vscale_core_DW01_inc_7_U255 ( .A1(vscale_core_DW01_inc_7n187), .A2(vscale_core_DW01_inc_7n180), .ZN(vscale_core_DW01_inc_7n179) );
  NOR2_X2 vscale_core_DW01_inc_7_U256 ( .A1(vscale_core_DW01_inc_7n132), .A2(vscale_core_DW01_inc_7n131), .ZN(vscale_core_DW01_inc_7n128) );
  NOR2_X2 vscale_core_DW01_inc_7_U257 ( .A1(vscale_core_DW01_inc_7n143), .A2(vscale_core_DW01_inc_7n142), .ZN(vscale_core_DW01_inc_7n139) );
  NOR2_X2 vscale_core_DW01_inc_7_U258 ( .A1(vscale_core_DW01_inc_7n153), .A2(vscale_core_DW01_inc_7n151), .ZN(vscale_core_DW01_inc_7n148) );
  NOR2_X2 vscale_core_DW01_inc_7_U259 ( .A1(vscale_core_DW01_inc_7n162), .A2(vscale_core_DW01_inc_7n161), .ZN(vscale_core_DW01_inc_7n158) );
  NOR2_X2 vscale_core_DW01_inc_7_U260 ( .A1(vscale_core_DW01_inc_7n187), .A2(vscale_core_DW01_inc_7n186), .ZN(vscale_core_DW01_inc_7n183) );
  NOR2_X2 vscale_core_DW01_inc_7_U261 ( .A1(vscale_core_DW01_inc_7n45), .A2(vscale_core_DW01_inc_7n43), .ZN(vscale_core_DW01_inc_7n40) );
  NOR2_X2 vscale_core_DW01_inc_7_U262 ( .A1(vscale_core_DW01_inc_7n54), .A2(vscale_core_DW01_inc_7n53), .ZN(vscale_core_DW01_inc_7n50) );
  NOR2_X2 vscale_core_DW01_inc_7_U263 ( .A1(vscale_core_DW01_inc_7n108), .A2(vscale_core_DW01_inc_7n101), .ZN(vscale_core_DW01_inc_7n100) );
  NOR2_X2 vscale_core_DW01_inc_7_U264 ( .A1(vscale_core_DW01_inc_7n180), .A2(vscale_core_DW01_inc_7n173), .ZN(vscale_core_DW01_inc_7n172) );
  NOR2_X2 vscale_core_DW01_inc_7_U265 ( .A1(vscale_core_DW01_inc_7n125), .A2(vscale_core_DW01_inc_7n118), .ZN(vscale_core_DW01_inc_7n117) );
  NOR2_X2 vscale_core_DW01_inc_7_U266 ( .A1(vscale_core_DW01_inc_7n189), .A2(vscale_core_DW01_inc_7n196), .ZN(vscale_core_DW01_inc_7n188) );
  NOR2_X2 vscale_core_DW01_inc_7_U267 ( .A1(vscale_core_DW01_inc_7n134), .A2(vscale_core_DW01_inc_7n171), .ZN(vscale_core_DW01_inc_7n133) );
  NOR2_X2 vscale_core_DW01_inc_7_U268 ( .A1(vscale_core_DW01_inc_7n145), .A2(vscale_core_DW01_inc_7n136), .ZN(vscale_core_DW01_inc_7n135) );
  NOR2_X2 vscale_core_DW01_inc_7_U269 ( .A1(vscale_core_DW01_inc_7n164), .A2(vscale_core_DW01_inc_7n155), .ZN(vscale_core_DW01_inc_7n154) );
  NOR2_X2 vscale_core_DW01_inc_7_U270 ( .A1(vscale_core_DW01_inc_7n63), .A2(vscale_core_DW01_inc_7n24), .ZN(vscale_core_DW01_inc_7n23) );
  NOR2_X2 vscale_core_DW01_inc_7_U271 ( .A1(vscale_core_DW01_inc_7n91), .A2(vscale_core_DW01_inc_7n84), .ZN(vscale_core_DW01_inc_7n83) );
  NOR2_X2 vscale_core_DW01_inc_7_U272 ( .A1(vscale_core_DW01_inc_7n56), .A2(vscale_core_DW01_inc_7n47), .ZN(vscale_core_DW01_inc_7n46) );
  INV_X4 vscale_core_DW01_inc_7_U273 ( .A(vscale_core_DW01_inc_7n98), .ZN(vscale_core_DW01_inc_7n97) );
  INV_X4 vscale_core_DW01_inc_7_U274 ( .A(pipeline_csr_cycle_full[24]), .ZN(vscale_core_DW01_inc_7n96) );
  INV_X4 vscale_core_DW01_inc_7_U275 ( .A(pipeline_csr_cycle_full[25]), .ZN(vscale_core_DW01_inc_7n93) );
  INV_X4 vscale_core_DW01_inc_7_U276 ( .A(pipeline_csr_cycle_full[26]), .ZN(vscale_core_DW01_inc_7n89) );
  INV_X4 vscale_core_DW01_inc_7_U277 ( .A(pipeline_csr_cycle_full[27]), .ZN(vscale_core_DW01_inc_7n86) );
  INV_X4 vscale_core_DW01_inc_7_U278 ( .A(vscale_core_DW01_inc_7n83), .ZN(vscale_core_DW01_inc_7n82) );
  INV_X4 vscale_core_DW01_inc_7_U279 ( .A(vscale_core_DW01_inc_7n81), .ZN(vscale_core_DW01_inc_7n80) );
  INV_X4 vscale_core_DW01_inc_7_U280 ( .A(pipeline_csr_cycle_full[28]), .ZN(vscale_core_DW01_inc_7n79) );
  INV_X4 vscale_core_DW01_inc_7_U281 ( .A(pipeline_csr_cycle_full[29]), .ZN(vscale_core_DW01_inc_7n76) );
  INV_X4 vscale_core_DW01_inc_7_U282 ( .A(pipeline_csr_cycle_full[30]), .ZN(vscale_core_DW01_inc_7n72) );
  INV_X4 vscale_core_DW01_inc_7_U283 ( .A(pipeline_csr_cycle_full[31]), .ZN(vscale_core_DW01_inc_7n69) );
  INV_X4 vscale_core_DW01_inc_7_U284 ( .A(vscale_core_DW01_inc_7n63), .ZN(vscale_core_DW01_inc_7n62) );
  INV_X4 vscale_core_DW01_inc_7_U285 ( .A(pipeline_csr_cycle_full[32]), .ZN(vscale_core_DW01_inc_7n61) );
  INV_X4 vscale_core_DW01_inc_7_U286 ( .A(pipeline_csr_cycle_full[33]), .ZN(vscale_core_DW01_inc_7n58) );
  INV_X4 vscale_core_DW01_inc_7_U287 ( .A(vscale_core_DW01_inc_7n56), .ZN(vscale_core_DW01_inc_7n55) );
  INV_X4 vscale_core_DW01_inc_7_U288 ( .A(pipeline_csr_cycle_full[34]), .ZN(vscale_core_DW01_inc_7n53) );
  INV_X4 vscale_core_DW01_inc_7_U289 ( .A(pipeline_csr_cycle_full[35]), .ZN(vscale_core_DW01_inc_7n49) );
  INV_X4 vscale_core_DW01_inc_7_U290 ( .A(vscale_core_DW01_inc_7n45), .ZN(vscale_core_DW01_inc_7n44) );
  INV_X4 vscale_core_DW01_inc_7_U291 ( .A(pipeline_csr_cycle_full[36]), .ZN(vscale_core_DW01_inc_7n43) );
  INV_X4 vscale_core_DW01_inc_7_U292 ( .A(pipeline_csr_cycle_full[37]), .ZN(vscale_core_DW01_inc_7n39) );
  INV_X4 vscale_core_DW01_inc_7_U293 ( .A(vscale_core_DW01_inc_7n37), .ZN(vscale_core_DW01_inc_7n36) );
  INV_X4 vscale_core_DW01_inc_7_U294 ( .A(pipeline_csr_cycle_full[38]), .ZN(vscale_core_DW01_inc_7n34) );
  INV_X4 vscale_core_DW01_inc_7_U295 ( .A(vscale_core_DW01_inc_7n32), .ZN(vscale_core_DW01_inc_7n31) );
  INV_X4 vscale_core_DW01_inc_7_U296 ( .A(pipeline_csr_cycle_full[39]), .ZN(vscale_core_DW01_inc_7n29) );
  INV_X4 vscale_core_DW01_inc_7_U297 ( .A(pipeline_csr_cycle_full[40]), .ZN(vscale_core_DW01_inc_7n26) );
  INV_X4 vscale_core_DW01_inc_7_U298 ( .A(pipeline_csr_cycle_full[1]), .ZN(vscale_core_DW01_inc_7n198) );
  INV_X4 vscale_core_DW01_inc_7_U299 ( .A(vscale_core_DW01_inc_7n196), .ZN(vscale_core_DW01_inc_7n195) );
  INV_X4 vscale_core_DW01_inc_7_U300 ( .A(pipeline_csr_cycle_full[2]), .ZN(vscale_core_DW01_inc_7n194) );
  INV_X4 vscale_core_DW01_inc_7_U301 ( .A(pipeline_csr_cycle_full[3]), .ZN(vscale_core_DW01_inc_7n191) );
  INV_X4 vscale_core_DW01_inc_7_U302 ( .A(vscale_core_DW01_inc_7n188), .ZN(vscale_core_DW01_inc_7n187) );
  INV_X4 vscale_core_DW01_inc_7_U303 ( .A(pipeline_csr_cycle_full[4]), .ZN(vscale_core_DW01_inc_7n186) );
  INV_X4 vscale_core_DW01_inc_7_U304 ( .A(pipeline_csr_cycle_full[5]), .ZN(vscale_core_DW01_inc_7n182) );
  INV_X4 vscale_core_DW01_inc_7_U305 ( .A(pipeline_csr_cycle_full[6]), .ZN(vscale_core_DW01_inc_7n178) );
  INV_X4 vscale_core_DW01_inc_7_U306 ( .A(pipeline_csr_cycle_full[7]), .ZN(vscale_core_DW01_inc_7n175) );
  INV_X4 vscale_core_DW01_inc_7_U307 ( .A(vscale_core_DW01_inc_7n171), .ZN(vscale_core_DW01_inc_7n170) );
  INV_X4 vscale_core_DW01_inc_7_U308 ( .A(pipeline_csr_cycle_full[8]), .ZN(vscale_core_DW01_inc_7n169) );
  INV_X4 vscale_core_DW01_inc_7_U309 ( .A(pipeline_csr_cycle_full[9]), .ZN(vscale_core_DW01_inc_7n166) );
  INV_X4 vscale_core_DW01_inc_7_U310 ( .A(vscale_core_DW01_inc_7n164), .ZN(vscale_core_DW01_inc_7n163) );
  INV_X4 vscale_core_DW01_inc_7_U311 ( .A(pipeline_csr_cycle_full[10]), .ZN(vscale_core_DW01_inc_7n161) );
  INV_X4 vscale_core_DW01_inc_7_U312 ( .A(pipeline_csr_cycle_full[11]), .ZN(vscale_core_DW01_inc_7n157) );
  INV_X4 vscale_core_DW01_inc_7_U313 ( .A(vscale_core_DW01_inc_7n153), .ZN(vscale_core_DW01_inc_7n152) );
  INV_X4 vscale_core_DW01_inc_7_U314 ( .A(pipeline_csr_cycle_full[12]), .ZN(vscale_core_DW01_inc_7n151) );
  INV_X4 vscale_core_DW01_inc_7_U315 ( .A(pipeline_csr_cycle_full[13]), .ZN(vscale_core_DW01_inc_7n147) );
  INV_X4 vscale_core_DW01_inc_7_U316 ( .A(vscale_core_DW01_inc_7n145), .ZN(vscale_core_DW01_inc_7n144) );
  INV_X4 vscale_core_DW01_inc_7_U317 ( .A(pipeline_csr_cycle_full[14]), .ZN(vscale_core_DW01_inc_7n142) );
  INV_X4 vscale_core_DW01_inc_7_U318 ( .A(pipeline_csr_cycle_full[15]), .ZN(vscale_core_DW01_inc_7n138) );
  INV_X4 vscale_core_DW01_inc_7_U319 ( .A(vscale_core_DW01_inc_7n133), .ZN(vscale_core_DW01_inc_7n132) );
  INV_X4 vscale_core_DW01_inc_7_U320 ( .A(pipeline_csr_cycle_full[16]), .ZN(vscale_core_DW01_inc_7n131) );
  INV_X4 vscale_core_DW01_inc_7_U321 ( .A(pipeline_csr_cycle_full[17]), .ZN(vscale_core_DW01_inc_7n127) );
  INV_X4 vscale_core_DW01_inc_7_U322 ( .A(pipeline_csr_cycle_full[18]), .ZN(vscale_core_DW01_inc_7n123) );
  INV_X4 vscale_core_DW01_inc_7_U323 ( .A(pipeline_csr_cycle_full[19]), .ZN(vscale_core_DW01_inc_7n120) );
  INV_X4 vscale_core_DW01_inc_7_U324 ( .A(vscale_core_DW01_inc_7n117), .ZN(vscale_core_DW01_inc_7n116) );
  INV_X4 vscale_core_DW01_inc_7_U325 ( .A(vscale_core_DW01_inc_7n115), .ZN(vscale_core_DW01_inc_7n114) );
  INV_X4 vscale_core_DW01_inc_7_U326 ( .A(pipeline_csr_cycle_full[20]), .ZN(vscale_core_DW01_inc_7n113) );
  INV_X4 vscale_core_DW01_inc_7_U327 ( .A(pipeline_csr_cycle_full[21]), .ZN(vscale_core_DW01_inc_7n110) );
  INV_X4 vscale_core_DW01_inc_7_U328 ( .A(pipeline_csr_cycle_full[22]), .ZN(vscale_core_DW01_inc_7n106) );
  INV_X4 vscale_core_DW01_inc_7_U329 ( .A(pipeline_csr_cycle_full[23]), .ZN(vscale_core_DW01_inc_7n103) );
  INV_X4 vscale_core_DW01_inc_7_U330 ( .A(pipeline_csr_cycle_full[0]), .ZN(pipeline_csr_N648) );
;
  vscale_core_DW01_add_8 pipeline_csr_add_218_aco 

  XOR2_X2 vscale_core_DW01_add_8_U1 ( .A(n12597), .B(vscale_core_DW01_add_8n3), .Z(pipeline_csr_N332) );
  HA_X1 vscale_core_DW01_add_8_U2 ( .A(n10794), .B(vscale_core_DW01_add_8n4), .CO(vscale_core_DW01_add_8n3), .S(pipeline_csr_N331) );
  HA_X1 vscale_core_DW01_add_8_U3 ( .A(n10795), .B(vscale_core_DW01_add_8n5), .CO(vscale_core_DW01_add_8n4), .S(pipeline_csr_N330) );
  HA_X1 vscale_core_DW01_add_8_U4 ( .A(n10796), .B(vscale_core_DW01_add_8n6), .CO(vscale_core_DW01_add_8n5), .S(pipeline_csr_N329) );
  HA_X1 vscale_core_DW01_add_8_U5 ( .A(n10797), .B(vscale_core_DW01_add_8n7), .CO(vscale_core_DW01_add_8n6), .S(pipeline_csr_N328) );
  HA_X1 vscale_core_DW01_add_8_U6 ( .A(n10799), .B(vscale_core_DW01_add_8n8), .CO(vscale_core_DW01_add_8n7), .S(pipeline_csr_N327) );
  HA_X1 vscale_core_DW01_add_8_U7 ( .A(n10800), .B(vscale_core_DW01_add_8n9), .CO(vscale_core_DW01_add_8n8), .S(pipeline_csr_N326) );
  HA_X1 vscale_core_DW01_add_8_U8 ( .A(n10801), .B(vscale_core_DW01_add_8n10), .CO(vscale_core_DW01_add_8n9), .S(pipeline_csr_N325) );
  HA_X1 vscale_core_DW01_add_8_U9 ( .A(n10802), .B(vscale_core_DW01_add_8n11), .CO(vscale_core_DW01_add_8n10), .S(pipeline_csr_N324) );
  HA_X1 vscale_core_DW01_add_8_U10 ( .A(n10803), .B(vscale_core_DW01_add_8n12), .CO(vscale_core_DW01_add_8n11), .S(pipeline_csr_N323) );
  HA_X1 vscale_core_DW01_add_8_U11 ( .A(n10804), .B(vscale_core_DW01_add_8n13), .CO(vscale_core_DW01_add_8n12), .S(pipeline_csr_N322) );
  HA_X1 vscale_core_DW01_add_8_U12 ( .A(n10805), .B(vscale_core_DW01_add_8n14), .CO(vscale_core_DW01_add_8n13), .S(pipeline_csr_N321) );
  HA_X1 vscale_core_DW01_add_8_U13 ( .A(n10806), .B(vscale_core_DW01_add_8n15), .CO(vscale_core_DW01_add_8n14), .S(pipeline_csr_N320) );
  HA_X1 vscale_core_DW01_add_8_U14 ( .A(n10807), .B(vscale_core_DW01_add_8n16), .CO(vscale_core_DW01_add_8n15), .S(pipeline_csr_N319) );
  HA_X1 vscale_core_DW01_add_8_U15 ( .A(n10809), .B(vscale_core_DW01_add_8n17), .CO(vscale_core_DW01_add_8n16), .S(pipeline_csr_N318) );
  HA_X1 vscale_core_DW01_add_8_U16 ( .A(n10810), .B(vscale_core_DW01_add_8n18), .CO(vscale_core_DW01_add_8n17), .S(pipeline_csr_N317) );
  HA_X1 vscale_core_DW01_add_8_U17 ( .A(n10811), .B(vscale_core_DW01_add_8n19), .CO(vscale_core_DW01_add_8n18), .S(pipeline_csr_N316) );
  HA_X1 vscale_core_DW01_add_8_U18 ( .A(n10812), .B(vscale_core_DW01_add_8n20), .CO(vscale_core_DW01_add_8n19), .S(pipeline_csr_N315) );
  HA_X1 vscale_core_DW01_add_8_U19 ( .A(n10813), .B(vscale_core_DW01_add_8n21), .CO(vscale_core_DW01_add_8n20), .S(pipeline_csr_N314) );
  HA_X1 vscale_core_DW01_add_8_U20 ( .A(n10814), .B(vscale_core_DW01_add_8n22), .CO(vscale_core_DW01_add_8n21), .S(pipeline_csr_N313) );
  HA_X1 vscale_core_DW01_add_8_U21 ( .A(n10815), .B(vscale_core_DW01_add_8n23), .CO(vscale_core_DW01_add_8n22), .S(pipeline_csr_N312) );
  HA_X1 vscale_core_DW01_add_8_U22 ( .A(n10816), .B(vscale_core_DW01_add_8n24), .CO(vscale_core_DW01_add_8n23), .S(pipeline_csr_N311) );
  HA_X1 vscale_core_DW01_add_8_U23 ( .A(n10817), .B(vscale_core_DW01_add_8n25), .CO(vscale_core_DW01_add_8n24), .S(pipeline_csr_N310) );
  HA_X1 vscale_core_DW01_add_8_U24 ( .A(n10818), .B(vscale_core_DW01_add_8n26), .CO(vscale_core_DW01_add_8n25), .S(pipeline_csr_N309) );
  HA_X1 vscale_core_DW01_add_8_U25 ( .A(n10819), .B(vscale_core_DW01_add_8n144), .CO(vscale_core_DW01_add_8n26), .S(pipeline_csr_N308) );
  XNOR2_X2 vscale_core_DW01_add_8_U27 ( .A(vscale_core_DW01_add_8n30), .B(vscale_core_DW01_add_8n29), .ZN(pipeline_csr_N307) );
  XOR2_X2 vscale_core_DW01_add_8_U31 ( .A(vscale_core_DW01_add_8n31), .B(vscale_core_DW01_add_8n32), .Z(pipeline_csr_N306) );
  XNOR2_X2 vscale_core_DW01_add_8_U34 ( .A(vscale_core_DW01_add_8n37), .B(vscale_core_DW01_add_8n36), .ZN(pipeline_csr_N305) );
  NAND2_X2 vscale_core_DW01_add_8_U37 ( .A1(n12144), .A2(n12808), .ZN(vscale_core_DW01_add_8n34) );
  XOR2_X2 vscale_core_DW01_add_8_U40 ( .A(vscale_core_DW01_add_8n40), .B(vscale_core_DW01_add_8n1), .Z(pipeline_csr_N304) );
  NAND2_X2 vscale_core_DW01_add_8_U49 ( .A1(n6369), .A2(n12290), .ZN(vscale_core_DW01_add_8n1) );
  AND2_X4 vscale_core_DW01_add_8_U53 ( .A1(vscale_core_DW01_add_8n33), .A2(vscale_core_DW01_add_8n28), .ZN(vscale_core_DW01_add_8n144) );
  AND2_X4 vscale_core_DW01_add_8_U54 ( .A1(vscale_core_DW01_add_8n146), .A2(vscale_core_DW01_add_8n1), .ZN(pipeline_csr_N303) );
  NOR2_X2 vscale_core_DW01_add_8_U55 ( .A1(vscale_core_DW01_add_8n1), .A2(vscale_core_DW01_add_8n40), .ZN(vscale_core_DW01_add_8n37) );
  NOR2_X2 vscale_core_DW01_add_8_U56 ( .A1(vscale_core_DW01_add_8n1), .A2(vscale_core_DW01_add_8n34), .ZN(vscale_core_DW01_add_8n33) );
  NOR2_X2 vscale_core_DW01_add_8_U57 ( .A1(vscale_core_DW01_add_8n31), .A2(vscale_core_DW01_add_8n29), .ZN(vscale_core_DW01_add_8n28) );
  NOR2_X2 vscale_core_DW01_add_8_U58 ( .A1(vscale_core_DW01_add_8n32), .A2(vscale_core_DW01_add_8n31), .ZN(vscale_core_DW01_add_8n30) );
  OR2_X1 vscale_core_DW01_add_8_U59 ( .A1(n6369), .A2(n12290), .ZN(vscale_core_DW01_add_8n146) );
  INV_X4 vscale_core_DW01_add_8_U60 ( .A(n12144), .ZN(vscale_core_DW01_add_8n40) );
  INV_X4 vscale_core_DW01_add_8_U61 ( .A(n12808), .ZN(vscale_core_DW01_add_8n36) );
  INV_X4 vscale_core_DW01_add_8_U62 ( .A(vscale_core_DW01_add_8n33), .ZN(vscale_core_DW01_add_8n32) );
  INV_X4 vscale_core_DW01_add_8_U63 ( .A(n10822), .ZN(vscale_core_DW01_add_8n31) );
  INV_X4 vscale_core_DW01_add_8_U64 ( .A(n10820), .ZN(vscale_core_DW01_add_8n29) );
;
  vscale_core_DW01_add_9 pipeline_csr_add_92 

  XOR2_X2 vscale_core_DW01_add_9_U1 ( .A(n10282), .B(vscale_core_DW01_add_9n4), .Z(pipeline_handler_PC[31]) );
  HA_X1 vscale_core_DW01_add_9_U2 ( .A(n10238), .B(vscale_core_DW01_add_9n5), .CO(vscale_core_DW01_add_9n4), .S(pipeline_handler_PC[30]) );
  HA_X1 vscale_core_DW01_add_9_U3 ( .A(n10358), .B(vscale_core_DW01_add_9n6), .CO(vscale_core_DW01_add_9n5), .S(pipeline_handler_PC[29]) );
  HA_X1 vscale_core_DW01_add_9_U4 ( .A(n10426), .B(vscale_core_DW01_add_9n7), .CO(vscale_core_DW01_add_9n6), .S(pipeline_handler_PC[28]) );
  HA_X1 vscale_core_DW01_add_9_U5 ( .A(n10461), .B(vscale_core_DW01_add_9n8), .CO(vscale_core_DW01_add_9n7), .S(pipeline_handler_PC[27]) );
  HA_X1 vscale_core_DW01_add_9_U6 ( .A(n10537), .B(vscale_core_DW01_add_9n9), .CO(vscale_core_DW01_add_9n8), .S(pipeline_handler_PC[26]) );
  HA_X1 vscale_core_DW01_add_9_U7 ( .A(n10591), .B(vscale_core_DW01_add_9n10), .CO(vscale_core_DW01_add_9n9), .S(pipeline_handler_PC[25]) );
  HA_X1 vscale_core_DW01_add_9_U8 ( .A(n10645), .B(vscale_core_DW01_add_9n11), .CO(vscale_core_DW01_add_9n10), .S(pipeline_handler_PC[24]) );
  HA_X1 vscale_core_DW01_add_9_U9 ( .A(n10699), .B(vscale_core_DW01_add_9n12), .CO(vscale_core_DW01_add_9n11), .S(pipeline_handler_PC[23]) );
  HA_X1 vscale_core_DW01_add_9_U10 ( .A(n10750), .B(vscale_core_DW01_add_9n13), .CO(vscale_core_DW01_add_9n12), .S(pipeline_handler_PC[22]) );
  HA_X1 vscale_core_DW01_add_9_U11 ( .A(n10835), .B(vscale_core_DW01_add_9n14), .CO(vscale_core_DW01_add_9n13), .S(pipeline_handler_PC[21]) );
  HA_X1 vscale_core_DW01_add_9_U12 ( .A(n10895), .B(vscale_core_DW01_add_9n15), .CO(vscale_core_DW01_add_9n14), .S(pipeline_handler_PC[20]) );
  HA_X1 vscale_core_DW01_add_9_U13 ( .A(n10943), .B(vscale_core_DW01_add_9n16), .CO(vscale_core_DW01_add_9n15), .S(pipeline_handler_PC[19]) );
  HA_X1 vscale_core_DW01_add_9_U14 ( .A(n11003), .B(vscale_core_DW01_add_9n17), .CO(vscale_core_DW01_add_9n16), .S(pipeline_handler_PC[18]) );
  HA_X1 vscale_core_DW01_add_9_U15 ( .A(n11050), .B(vscale_core_DW01_add_9n18), .CO(vscale_core_DW01_add_9n17), .S(pipeline_handler_PC[17]) );
  HA_X1 vscale_core_DW01_add_9_U16 ( .A(n11077), .B(vscale_core_DW01_add_9n19), .CO(vscale_core_DW01_add_9n18), .S(pipeline_handler_PC[16]) );
  HA_X1 vscale_core_DW01_add_9_U17 ( .A(n11113), .B(vscale_core_DW01_add_9n20), .CO(vscale_core_DW01_add_9n19), .S(pipeline_handler_PC[15]) );
  HA_X1 vscale_core_DW01_add_9_U18 ( .A(n11133), .B(vscale_core_DW01_add_9n21), .CO(vscale_core_DW01_add_9n20), .S(pipeline_handler_PC[14]) );
  HA_X1 vscale_core_DW01_add_9_U19 ( .A(n11023), .B(vscale_core_DW01_add_9n22), .CO(vscale_core_DW01_add_9n21), .S(pipeline_handler_PC[13]) );
  HA_X1 vscale_core_DW01_add_9_U20 ( .A(n10862), .B(vscale_core_DW01_add_9n23), .CO(vscale_core_DW01_add_9n22), .S(pipeline_handler_PC[12]) );
  HA_X1 vscale_core_DW01_add_9_U21 ( .A(n10916), .B(vscale_core_DW01_add_9n24), .CO(vscale_core_DW01_add_9n23), .S(pipeline_handler_PC[11]) );
  HA_X1 vscale_core_DW01_add_9_U22 ( .A(n10970), .B(vscale_core_DW01_add_9n139), .CO(vscale_core_DW01_add_9n24), .S(pipeline_handler_PC[10]) );
  XNOR2_X2 vscale_core_DW01_add_9_U24 ( .A(vscale_core_DW01_add_9n28), .B(vscale_core_DW01_add_9n27), .ZN(pipeline_handler_PC[9]) );
  XNOR2_X2 vscale_core_DW01_add_9_U28 ( .A(vscale_core_DW01_add_9n32), .B(vscale_core_DW01_add_9n31), .ZN(pipeline_handler_PC[8]) );
  NAND2_X2 vscale_core_DW01_add_9_U31 ( .A1(n10673), .A2(n10635), .ZN(vscale_core_DW01_add_9n29) );
  XNOR2_X2 vscale_core_DW01_add_9_U34 ( .A(vscale_core_DW01_add_9n36), .B(vscale_core_DW01_add_9n35), .ZN(pipeline_handler_PC[7]) );
  FA_X1 vscale_core_DW01_add_9_U40 ( .A(pipeline_ctrl_N82), .B(pipeline_csr_mtvec[6]), .CI(vscale_core_DW01_add_9n40), .CO(vscale_core_DW01_add_9n36), .S(pipeline_handler_PC[6]) );
  NAND2_X2 vscale_core_DW01_add_9_U46 ( .A1(pipeline_csr_mtvec[5]), .A2(pipeline_ctrl_N81), .ZN(vscale_core_DW01_add_9n38) );
  AND2_X4 vscale_core_DW01_add_9_U50 ( .A1(vscale_core_DW01_add_9n36), .A2(vscale_core_DW01_add_9n26), .ZN(vscale_core_DW01_add_9n139) );
  AND2_X4 vscale_core_DW01_add_9_U51 ( .A1(vscale_core_DW01_add_9n141), .A2(vscale_core_DW01_add_9n38), .ZN(pipeline_handler_PC[5]) );
  INV_X1 vscale_core_DW01_add_9_U52 ( .A(vscale_core_DW01_add_9n36), .ZN(vscale_core_DW01_add_9n2) );
  NOR2_X2 vscale_core_DW01_add_9_U53 ( .A1(vscale_core_DW01_add_9n2), .A2(vscale_core_DW01_add_9n29), .ZN(vscale_core_DW01_add_9n28) );
  NOR2_X2 vscale_core_DW01_add_9_U54 ( .A1(vscale_core_DW01_add_9n2), .A2(vscale_core_DW01_add_9n35), .ZN(vscale_core_DW01_add_9n32) );
  NOR2_X2 vscale_core_DW01_add_9_U55 ( .A1(vscale_core_DW01_add_9n29), .A2(vscale_core_DW01_add_9n27), .ZN(vscale_core_DW01_add_9n26) );
  OR2_X1 vscale_core_DW01_add_9_U56 ( .A1(pipeline_csr_mtvec[5]), .A2(pipeline_ctrl_N81), .ZN(vscale_core_DW01_add_9n141) );
  BUF_X4 vscale_core_DW01_add_9_U57 ( .A(pipeline_csr_mtvec[2]), .Z(pipeline_handler_PC[2]) );
  BUF_X4 vscale_core_DW01_add_9_U58 ( .A(pipeline_csr_mtvec[3]), .Z(pipeline_handler_PC[3]) );
  BUF_X4 vscale_core_DW01_add_9_U59 ( .A(pipeline_csr_mtvec[4]), .Z(pipeline_handler_PC[4]) );
  INV_X4 vscale_core_DW01_add_9_U60 ( .A(vscale_core_DW01_add_9n38), .ZN(vscale_core_DW01_add_9n40) );
  INV_X4 vscale_core_DW01_add_9_U61 ( .A(n10673), .ZN(vscale_core_DW01_add_9n35) );
  INV_X4 vscale_core_DW01_add_9_U62 ( .A(n10635), .ZN(vscale_core_DW01_add_9n31) );
  INV_X4 vscale_core_DW01_add_9_U63 ( .A(n10564), .ZN(vscale_core_DW01_add_9n27) );
;
  vscale_core_DW01_add_10 pipeline_PCmux_add_55 

  XNOR2_X2 vscale_core_DW01_add_10_U5 ( .A(vscale_core_DW01_add_10n38), .B(vscale_core_DW01_add_10n5), .ZN(n13160) );
  NAND2_X2 vscale_core_DW01_add_10_U6 ( .A1(vscale_core_DW01_add_10n406), .A2(vscale_core_DW01_add_10n37), .ZN(vscale_core_DW01_add_10n5) );
  NAND2_X2 vscale_core_DW01_add_10_U9 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[31]), .ZN(vscale_core_DW01_add_10n37) );
  XNOR2_X2 vscale_core_DW01_add_10_U10 ( .A(vscale_core_DW01_add_10n49), .B(vscale_core_DW01_add_10n6), .ZN(n13161) );
  NAND2_X2 vscale_core_DW01_add_10_U20 ( .A1(vscale_core_DW01_add_10n279), .A2(vscale_core_DW01_add_10n48), .ZN(vscale_core_DW01_add_10n6) );
  XNOR2_X2 vscale_core_DW01_add_10_U24 ( .A(vscale_core_DW01_add_10n58), .B(vscale_core_DW01_add_10n7), .ZN(n13162) );
  NAND2_X2 vscale_core_DW01_add_10_U32 ( .A1(vscale_core_DW01_add_10n280), .A2(vscale_core_DW01_add_10n57), .ZN(vscale_core_DW01_add_10n7) );
  NAND2_X2 vscale_core_DW01_add_10_U35 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[29]), .ZN(vscale_core_DW01_add_10n57) );
  XNOR2_X2 vscale_core_DW01_add_10_U36 ( .A(vscale_core_DW01_add_10n69), .B(vscale_core_DW01_add_10n8), .ZN(n13163) );
  NAND2_X2 vscale_core_DW01_add_10_U42 ( .A1(vscale_core_DW01_add_10n81), .A2(vscale_core_DW01_add_10n65), .ZN(vscale_core_DW01_add_10n63) );
  NAND2_X2 vscale_core_DW01_add_10_U46 ( .A1(vscale_core_DW01_add_10n281), .A2(vscale_core_DW01_add_10n68), .ZN(vscale_core_DW01_add_10n8) );
  XNOR2_X2 vscale_core_DW01_add_10_U50 ( .A(vscale_core_DW01_add_10n78), .B(vscale_core_DW01_add_10n9), .ZN(n13164) );
  NAND2_X2 vscale_core_DW01_add_10_U58 ( .A1(vscale_core_DW01_add_10n282), .A2(vscale_core_DW01_add_10n77), .ZN(vscale_core_DW01_add_10n9) );
  NAND2_X2 vscale_core_DW01_add_10_U61 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[27]), .ZN(vscale_core_DW01_add_10n77) );
  XNOR2_X2 vscale_core_DW01_add_10_U62 ( .A(vscale_core_DW01_add_10n89), .B(vscale_core_DW01_add_10n10), .ZN(n13165) );
  NAND2_X2 vscale_core_DW01_add_10_U72 ( .A1(vscale_core_DW01_add_10n283), .A2(vscale_core_DW01_add_10n88), .ZN(vscale_core_DW01_add_10n10) );
  NAND2_X2 vscale_core_DW01_add_10_U75 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[26]), .ZN(vscale_core_DW01_add_10n88) );
  XNOR2_X2 vscale_core_DW01_add_10_U76 ( .A(vscale_core_DW01_add_10n96), .B(vscale_core_DW01_add_10n11), .ZN(n13166) );
  NAND2_X2 vscale_core_DW01_add_10_U82 ( .A1(vscale_core_DW01_add_10n92), .A2(vscale_core_DW01_add_10n95), .ZN(vscale_core_DW01_add_10n11) );
  XNOR2_X2 vscale_core_DW01_add_10_U86 ( .A(vscale_core_DW01_add_10n107), .B(vscale_core_DW01_add_10n12), .ZN(n13167) );
  NAND2_X2 vscale_core_DW01_add_10_U92 ( .A1(vscale_core_DW01_add_10n119), .A2(vscale_core_DW01_add_10n103), .ZN(vscale_core_DW01_add_10n101) );
  NAND2_X2 vscale_core_DW01_add_10_U96 ( .A1(vscale_core_DW01_add_10n285), .A2(vscale_core_DW01_add_10n106), .ZN(vscale_core_DW01_add_10n12) );
  XNOR2_X2 vscale_core_DW01_add_10_U100 ( .A(vscale_core_DW01_add_10n116), .B(vscale_core_DW01_add_10n13), .ZN(n13168) );
  NAND2_X2 vscale_core_DW01_add_10_U102 ( .A1(vscale_core_DW01_add_10n110), .A2(vscale_core_DW01_add_10n137), .ZN(vscale_core_DW01_add_10n108) );
  NAND2_X2 vscale_core_DW01_add_10_U108 ( .A1(vscale_core_DW01_add_10n286), .A2(vscale_core_DW01_add_10n115), .ZN(vscale_core_DW01_add_10n13) );
  NAND2_X2 vscale_core_DW01_add_10_U111 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[23]), .ZN(vscale_core_DW01_add_10n115) );
  XNOR2_X2 vscale_core_DW01_add_10_U112 ( .A(vscale_core_DW01_add_10n127), .B(vscale_core_DW01_add_10n14), .ZN(n13169) );
  NAND2_X2 vscale_core_DW01_add_10_U114 ( .A1(vscale_core_DW01_add_10n137), .A2(vscale_core_DW01_add_10n119), .ZN(vscale_core_DW01_add_10n117) );
  NAND2_X2 vscale_core_DW01_add_10_U122 ( .A1(vscale_core_DW01_add_10n287), .A2(vscale_core_DW01_add_10n126), .ZN(vscale_core_DW01_add_10n14) );
  NAND2_X2 vscale_core_DW01_add_10_U125 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[22]), .ZN(vscale_core_DW01_add_10n126) );
  XNOR2_X2 vscale_core_DW01_add_10_U126 ( .A(vscale_core_DW01_add_10n134), .B(vscale_core_DW01_add_10n15), .ZN(n13170) );
  NAND2_X2 vscale_core_DW01_add_10_U128 ( .A1(vscale_core_DW01_add_10n137), .A2(vscale_core_DW01_add_10n288), .ZN(vscale_core_DW01_add_10n128) );
  NAND2_X2 vscale_core_DW01_add_10_U132 ( .A1(vscale_core_DW01_add_10n288), .A2(vscale_core_DW01_add_10n133), .ZN(vscale_core_DW01_add_10n15) );
  NAND2_X2 vscale_core_DW01_add_10_U135 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[21]), .ZN(vscale_core_DW01_add_10n133) );
  XNOR2_X2 vscale_core_DW01_add_10_U136 ( .A(vscale_core_DW01_add_10n145), .B(vscale_core_DW01_add_10n16), .ZN(n13171) );
  NAND2_X2 vscale_core_DW01_add_10_U142 ( .A1(vscale_core_DW01_add_10n141), .A2(vscale_core_DW01_add_10n155), .ZN(vscale_core_DW01_add_10n135) );
  AOI21_X4 vscale_core_DW01_add_10_U143 ( .B1(vscale_core_DW01_add_10n141), .B2(vscale_core_DW01_add_10n156), .A(vscale_core_DW01_add_10n142), .ZN(vscale_core_DW01_add_10n136) );
  NAND2_X2 vscale_core_DW01_add_10_U146 ( .A1(vscale_core_DW01_add_10n289), .A2(vscale_core_DW01_add_10n144), .ZN(vscale_core_DW01_add_10n16) );
  NAND2_X2 vscale_core_DW01_add_10_U149 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[20]), .ZN(vscale_core_DW01_add_10n144) );
  XNOR2_X2 vscale_core_DW01_add_10_U150 ( .A(vscale_core_DW01_add_10n152), .B(vscale_core_DW01_add_10n17), .ZN(n13172) );
  NAND2_X2 vscale_core_DW01_add_10_U152 ( .A1(vscale_core_DW01_add_10n155), .A2(vscale_core_DW01_add_10n290), .ZN(vscale_core_DW01_add_10n146) );
  NAND2_X2 vscale_core_DW01_add_10_U156 ( .A1(vscale_core_DW01_add_10n290), .A2(vscale_core_DW01_add_10n151), .ZN(vscale_core_DW01_add_10n17) );
  XNOR2_X2 vscale_core_DW01_add_10_U160 ( .A(vscale_core_DW01_add_10n163), .B(vscale_core_DW01_add_10n18), .ZN(n13173) );
  OAI21_X4 vscale_core_DW01_add_10_U169 ( .B1(vscale_core_DW01_add_10n161), .B2(vscale_core_DW01_add_10n165), .A(vscale_core_DW01_add_10n162), .ZN(vscale_core_DW01_add_10n156) );
  NAND2_X2 vscale_core_DW01_add_10_U170 ( .A1(vscale_core_DW01_add_10n291), .A2(vscale_core_DW01_add_10n162), .ZN(vscale_core_DW01_add_10n18) );
  XNOR2_X2 vscale_core_DW01_add_10_U180 ( .A(vscale_core_DW01_add_10n175), .B(vscale_core_DW01_add_10n20), .ZN(n13175) );
  NAND2_X2 vscale_core_DW01_add_10_U184 ( .A1(vscale_core_DW01_add_10n187), .A2(vscale_core_DW01_add_10n171), .ZN(vscale_core_DW01_add_10n169) );
  XNOR2_X2 vscale_core_DW01_add_10_U192 ( .A(vscale_core_DW01_add_10n184), .B(vscale_core_DW01_add_10n21), .ZN(n13176) );
  NAND2_X2 vscale_core_DW01_add_10_U194 ( .A1(vscale_core_DW01_add_10n178), .A2(vscale_core_DW01_add_10n205), .ZN(vscale_core_DW01_add_10n176) );
  XNOR2_X2 vscale_core_DW01_add_10_U204 ( .A(vscale_core_DW01_add_10n195), .B(vscale_core_DW01_add_10n22), .ZN(n13177) );
  NAND2_X2 vscale_core_DW01_add_10_U206 ( .A1(vscale_core_DW01_add_10n205), .A2(vscale_core_DW01_add_10n187), .ZN(vscale_core_DW01_add_10n185) );
  NAND2_X2 vscale_core_DW01_add_10_U214 ( .A1(vscale_core_DW01_add_10n295), .A2(vscale_core_DW01_add_10n194), .ZN(vscale_core_DW01_add_10n22) );
  XNOR2_X2 vscale_core_DW01_add_10_U218 ( .A(vscale_core_DW01_add_10n202), .B(vscale_core_DW01_add_10n23), .ZN(n13178) );
  NAND2_X2 vscale_core_DW01_add_10_U220 ( .A1(vscale_core_DW01_add_10n205), .A2(vscale_core_DW01_add_10n296), .ZN(vscale_core_DW01_add_10n196) );
  XNOR2_X2 vscale_core_DW01_add_10_U228 ( .A(vscale_core_DW01_add_10n213), .B(vscale_core_DW01_add_10n24), .ZN(n13179) );
  NAND2_X2 vscale_core_DW01_add_10_U241 ( .A1(pipeline_PCmux_base[12]), .A2(pipeline_PCmux_offset[12]), .ZN(vscale_core_DW01_add_10n212) );
  XNOR2_X2 vscale_core_DW01_add_10_U242 ( .A(vscale_core_DW01_add_10n220), .B(vscale_core_DW01_add_10n25), .ZN(n13180) );
  XNOR2_X2 vscale_core_DW01_add_10_U252 ( .A(vscale_core_DW01_add_10n231), .B(vscale_core_DW01_add_10n26), .ZN(n13181) );
  NAND2_X2 vscale_core_DW01_add_10_U265 ( .A1(pipeline_PCmux_base[10]), .A2(pipeline_PCmux_offset[10]), .ZN(vscale_core_DW01_add_10n230) );
  NAND2_X2 vscale_core_DW01_add_10_U271 ( .A1(pipeline_PCmux_base[9]), .A2(pipeline_PCmux_offset[9]), .ZN(vscale_core_DW01_add_10n233) );
  XOR2_X2 vscale_core_DW01_add_10_U272 ( .A(vscale_core_DW01_add_10n28), .B(vscale_core_DW01_add_10n242), .Z(n13183) );
  NAND2_X2 vscale_core_DW01_add_10_U275 ( .A1(vscale_core_DW01_add_10n250), .A2(vscale_core_DW01_add_10n238), .ZN(vscale_core_DW01_add_10n236) );
  NAND2_X2 vscale_core_DW01_add_10_U282 ( .A1(pipeline_PCmux_base[8]), .A2(pipeline_PCmux_offset[8]), .ZN(vscale_core_DW01_add_10n241) );
  XOR2_X2 vscale_core_DW01_add_10_U283 ( .A(vscale_core_DW01_add_10n29), .B(vscale_core_DW01_add_10n249), .Z(n13184) );
  NAND2_X2 vscale_core_DW01_add_10_U292 ( .A1(pipeline_PCmux_base[7]), .A2(pipeline_PCmux_offset[7]), .ZN(vscale_core_DW01_add_10n248) );
  XOR2_X2 vscale_core_DW01_add_10_U293 ( .A(vscale_core_DW01_add_10n30), .B(vscale_core_DW01_add_10n258), .Z(n13185) );
  NAND2_X2 vscale_core_DW01_add_10_U301 ( .A1(vscale_core_DW01_add_10n303), .A2(vscale_core_DW01_add_10n257), .ZN(vscale_core_DW01_add_10n30) );
  NAND2_X2 vscale_core_DW01_add_10_U304 ( .A1(pipeline_PCmux_base[6]), .A2(pipeline_PCmux_offset[6]), .ZN(vscale_core_DW01_add_10n257) );
  XNOR2_X2 vscale_core_DW01_add_10_U305 ( .A(vscale_core_DW01_add_10n263), .B(vscale_core_DW01_add_10n31), .ZN(imem_haddr[5]) );
  NAND2_X2 vscale_core_DW01_add_10_U309 ( .A1(vscale_core_DW01_add_10n304), .A2(vscale_core_DW01_add_10n262), .ZN(vscale_core_DW01_add_10n31) );
  XNOR2_X2 vscale_core_DW01_add_10_U313 ( .A(vscale_core_DW01_add_10n269), .B(vscale_core_DW01_add_10n32), .ZN(imem_haddr[4]) );
  NAND2_X2 vscale_core_DW01_add_10_U318 ( .A1(vscale_core_DW01_add_10n305), .A2(vscale_core_DW01_add_10n268), .ZN(vscale_core_DW01_add_10n32) );
  XOR2_X2 vscale_core_DW01_add_10_U328 ( .A(vscale_core_DW01_add_10n277), .B(vscale_core_DW01_add_10n34), .Z(imem_haddr[2]) );
  NAND2_X2 vscale_core_DW01_add_10_U331 ( .A1(vscale_core_DW01_add_10n307), .A2(vscale_core_DW01_add_10n275), .ZN(vscale_core_DW01_add_10n34) );
  NAND2_X2 vscale_core_DW01_add_10_U334 ( .A1(pipeline_PCmux_base[2]), .A2(pipeline_PCmux_offset[2]), .ZN(vscale_core_DW01_add_10n275) );
  NAND2_X2 vscale_core_DW01_add_10_U339 ( .A1(pipeline_PCmux_base[1]), .A2(pipeline_PCmux_offset[1]), .ZN(vscale_core_DW01_add_10n277) );
  AOI21_X2 vscale_core_DW01_add_10_U343 ( .B1(vscale_core_DW01_add_10n171), .B2(vscale_core_DW01_add_10n188), .A(vscale_core_DW01_add_10n172), .ZN(vscale_core_DW01_add_10n170) );
  OAI21_X1 vscale_core_DW01_add_10_U344 ( .B1(vscale_core_DW01_add_10n211), .B2(vscale_core_DW01_add_10n219), .A(vscale_core_DW01_add_10n212), .ZN(vscale_core_DW01_add_10n210) );
  NOR2_X4 vscale_core_DW01_add_10_U345 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[28]), .ZN(vscale_core_DW01_add_10n67) );
  AOI21_X4 vscale_core_DW01_add_10_U346 ( .B1(vscale_core_DW01_add_10n3), .B2(vscale_core_DW01_add_10n52), .A(vscale_core_DW01_add_10n53), .ZN(vscale_core_DW01_add_10n51) );
  AOI21_X4 vscale_core_DW01_add_10_U347 ( .B1(vscale_core_DW01_add_10n3), .B2(vscale_core_DW01_add_10n41), .A(vscale_core_DW01_add_10n42), .ZN(vscale_core_DW01_add_10n40) );
  OAI21_X4 vscale_core_DW01_add_10_U348 ( .B1(vscale_core_DW01_add_10n136), .B2(vscale_core_DW01_add_10n101), .A(vscale_core_DW01_add_10n102), .ZN(vscale_core_DW01_add_10n3) );
  NOR2_X4 vscale_core_DW01_add_10_U349 ( .A1(vscale_core_DW01_add_10n180), .A2(vscale_core_DW01_add_10n173), .ZN(vscale_core_DW01_add_10n171) );
  OAI21_X4 vscale_core_DW01_add_10_U350 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n164), .A(vscale_core_DW01_add_10n165), .ZN(vscale_core_DW01_add_10n163) );
  INV_X16 vscale_core_DW01_add_10_U351 ( .A(vscale_core_DW01_add_10n408), .ZN(vscale_core_DW01_add_10n409) );
  INV_X1 vscale_core_DW01_add_10_U352 ( .A(vscale_core_DW01_add_10n273), .ZN(vscale_core_DW01_add_10n272) );
  NOR2_X2 vscale_core_DW01_add_10_U353 ( .A1(vscale_core_DW01_add_10n203), .A2(vscale_core_DW01_add_10n169), .ZN(vscale_core_DW01_add_10n167) );
  NAND2_X1 vscale_core_DW01_add_10_U354 ( .A1(vscale_core_DW01_add_10n223), .A2(vscale_core_DW01_add_10n209), .ZN(vscale_core_DW01_add_10n203) );
  AOI21_X4 vscale_core_DW01_add_10_U355 ( .B1(vscale_core_DW01_add_10n235), .B2(vscale_core_DW01_add_10n167), .A(vscale_core_DW01_add_10n168), .ZN(vscale_core_DW01_add_10n2) );
  NOR2_X4 vscale_core_DW01_add_10_U356 ( .A1(pipeline_PCmux_base[8]), .A2(pipeline_PCmux_offset[8]), .ZN(vscale_core_DW01_add_10n240) );
  AOI21_X4 vscale_core_DW01_add_10_U357 ( .B1(vscale_core_DW01_add_10n65), .B2(vscale_core_DW01_add_10n82), .A(vscale_core_DW01_add_10n66), .ZN(vscale_core_DW01_add_10n64) );
  NOR2_X2 vscale_core_DW01_add_10_U358 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[22]), .ZN(vscale_core_DW01_add_10n125) );
  NOR2_X2 vscale_core_DW01_add_10_U359 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[24]), .ZN(vscale_core_DW01_add_10n105) );
  NOR2_X2 vscale_core_DW01_add_10_U360 ( .A1(pipeline_PCmux_base[6]), .A2(pipeline_PCmux_offset[6]), .ZN(vscale_core_DW01_add_10n256) );
  OAI21_X2 vscale_core_DW01_add_10_U361 ( .B1(vscale_core_DW01_add_10n193), .B2(vscale_core_DW01_add_10n201), .A(vscale_core_DW01_add_10n194), .ZN(vscale_core_DW01_add_10n188) );
  OAI21_X2 vscale_core_DW01_add_10_U362 ( .B1(vscale_core_DW01_add_10n256), .B2(vscale_core_DW01_add_10n262), .A(vscale_core_DW01_add_10n257), .ZN(vscale_core_DW01_add_10n251) );
  NOR2_X2 vscale_core_DW01_add_10_U363 ( .A1(vscale_core_DW01_add_10n261), .A2(vscale_core_DW01_add_10n256), .ZN(vscale_core_DW01_add_10n250) );
  NAND2_X2 vscale_core_DW01_add_10_U364 ( .A1(pipeline_PCmux_base[15]), .A2(pipeline_PCmux_offset[15]), .ZN(vscale_core_DW01_add_10n183) );
  INV_X4 vscale_core_DW01_add_10_U365 ( .A(vscale_core_DW01_add_10n2), .ZN(vscale_core_DW01_add_10n408) );
  NAND2_X2 vscale_core_DW01_add_10_U366 ( .A1(pipeline_PCmux_base[17]), .A2(pipeline_PCmux_offset[17]), .ZN(vscale_core_DW01_add_10n165) );
  AOI21_X2 vscale_core_DW01_add_10_U367 ( .B1(vscale_core_DW01_add_10n209), .B2(vscale_core_DW01_add_10n224), .A(vscale_core_DW01_add_10n210), .ZN(vscale_core_DW01_add_10n204) );
  NOR2_X2 vscale_core_DW01_add_10_U368 ( .A1(pipeline_PCmux_base[4]), .A2(pipeline_PCmux_offset[4]), .ZN(vscale_core_DW01_add_10n267) );
  NAND2_X2 vscale_core_DW01_add_10_U369 ( .A1(pipeline_PCmux_base[4]), .A2(pipeline_PCmux_offset[4]), .ZN(vscale_core_DW01_add_10n268) );
  OAI21_X2 vscale_core_DW01_add_10_U370 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n108), .A(vscale_core_DW01_add_10n109), .ZN(vscale_core_DW01_add_10n107) );
  OAI21_X2 vscale_core_DW01_add_10_U371 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n128), .A(vscale_core_DW01_add_10n129), .ZN(vscale_core_DW01_add_10n127) );
  OAI21_X2 vscale_core_DW01_add_10_U372 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n153), .A(vscale_core_DW01_add_10n154), .ZN(vscale_core_DW01_add_10n152) );
  OAI21_X2 vscale_core_DW01_add_10_U373 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n146), .A(vscale_core_DW01_add_10n147), .ZN(vscale_core_DW01_add_10n145) );
  NAND2_X1 vscale_core_DW01_add_10_U374 ( .A1(pipeline_PCmux_base[14]), .A2(pipeline_PCmux_offset[14]), .ZN(vscale_core_DW01_add_10n194) );
  NAND2_X1 vscale_core_DW01_add_10_U375 ( .A1(pipeline_PCmux_base[18]), .A2(pipeline_PCmux_offset[18]), .ZN(vscale_core_DW01_add_10n162) );
  NAND2_X2 vscale_core_DW01_add_10_U376 ( .A1(pipeline_PCmux_base[5]), .A2(pipeline_PCmux_offset[5]), .ZN(vscale_core_DW01_add_10n262) );
  NOR2_X1 vscale_core_DW01_add_10_U377 ( .A1(pipeline_PCmux_base[5]), .A2(pipeline_PCmux_offset[5]), .ZN(vscale_core_DW01_add_10n261) );
  AOI21_X2 vscale_core_DW01_add_10_U378 ( .B1(vscale_core_DW01_add_10n138), .B2(vscale_core_DW01_add_10n110), .A(vscale_core_DW01_add_10n111), .ZN(vscale_core_DW01_add_10n109) );
  NOR2_X2 vscale_core_DW01_add_10_U379 ( .A1(vscale_core_DW01_add_10n200), .A2(vscale_core_DW01_add_10n193), .ZN(vscale_core_DW01_add_10n187) );
  INV_X1 vscale_core_DW01_add_10_U380 ( .A(vscale_core_DW01_add_10n256), .ZN(vscale_core_DW01_add_10n303) );
  NOR2_X4 vscale_core_DW01_add_10_U381 ( .A1(pipeline_PCmux_base[10]), .A2(pipeline_PCmux_offset[10]), .ZN(vscale_core_DW01_add_10n229) );
  NOR2_X2 vscale_core_DW01_add_10_U382 ( .A1(vscale_core_DW01_add_10n132), .A2(vscale_core_DW01_add_10n125), .ZN(vscale_core_DW01_add_10n119) );
  OAI21_X2 vscale_core_DW01_add_10_U383 ( .B1(vscale_core_DW01_add_10n264), .B2(vscale_core_DW01_add_10n236), .A(vscale_core_DW01_add_10n237), .ZN(vscale_core_DW01_add_10n235) );
  OAI21_X2 vscale_core_DW01_add_10_U384 ( .B1(vscale_core_DW01_add_10n274), .B2(vscale_core_DW01_add_10n277), .A(vscale_core_DW01_add_10n275), .ZN(vscale_core_DW01_add_10n273) );
  NOR2_X2 vscale_core_DW01_add_10_U385 ( .A1(vscale_core_DW01_add_10n112), .A2(vscale_core_DW01_add_10n105), .ZN(vscale_core_DW01_add_10n103) );
  NOR2_X2 vscale_core_DW01_add_10_U386 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[20]), .ZN(vscale_core_DW01_add_10n143) );
  NOR2_X2 vscale_core_DW01_add_10_U387 ( .A1(pipeline_PCmux_base[18]), .A2(pipeline_PCmux_offset[18]), .ZN(vscale_core_DW01_add_10n161) );
  NOR2_X2 vscale_core_DW01_add_10_U388 ( .A1(pipeline_PCmux_base[14]), .A2(pipeline_PCmux_offset[14]), .ZN(vscale_core_DW01_add_10n193) );
  OAI21_X2 vscale_core_DW01_add_10_U389 ( .B1(vscale_core_DW01_add_10n229), .B2(vscale_core_DW01_add_10n233), .A(vscale_core_DW01_add_10n230), .ZN(vscale_core_DW01_add_10n224) );
  NOR2_X2 vscale_core_DW01_add_10_U390 ( .A1(pipeline_PCmux_base[12]), .A2(pipeline_PCmux_offset[12]), .ZN(vscale_core_DW01_add_10n211) );
  AOI21_X2 vscale_core_DW01_add_10_U391 ( .B1(vscale_core_DW01_add_10n273), .B2(vscale_core_DW01_add_10n265), .A(vscale_core_DW01_add_10n266), .ZN(vscale_core_DW01_add_10n264) );
  AOI21_X2 vscale_core_DW01_add_10_U392 ( .B1(vscale_core_DW01_add_10n138), .B2(vscale_core_DW01_add_10n288), .A(vscale_core_DW01_add_10n131), .ZN(vscale_core_DW01_add_10n129) );
  NOR2_X2 vscale_core_DW01_add_10_U393 ( .A1(pipeline_PCmux_base[17]), .A2(pipeline_PCmux_offset[17]), .ZN(vscale_core_DW01_add_10n164) );
  NAND2_X2 vscale_core_DW01_add_10_U394 ( .A1(pipeline_PCmux_base[13]), .A2(pipeline_PCmux_offset[13]), .ZN(vscale_core_DW01_add_10n201) );
  NOR2_X2 vscale_core_DW01_add_10_U395 ( .A1(pipeline_PCmux_base[2]), .A2(pipeline_PCmux_offset[2]), .ZN(vscale_core_DW01_add_10n274) );
  NAND2_X2 vscale_core_DW01_add_10_U396 ( .A1(pipeline_PCmux_base[3]), .A2(pipeline_PCmux_offset[3]), .ZN(vscale_core_DW01_add_10n271) );
  OAI21_X2 vscale_core_DW01_add_10_U397 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n97), .A(vscale_core_DW01_add_10n98), .ZN(vscale_core_DW01_add_10n96) );
  OAI21_X2 vscale_core_DW01_add_10_U398 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n135), .A(vscale_core_DW01_add_10n136), .ZN(vscale_core_DW01_add_10n134) );
  AOI21_X2 vscale_core_DW01_add_10_U399 ( .B1(vscale_core_DW01_add_10n103), .B2(vscale_core_DW01_add_10n120), .A(vscale_core_DW01_add_10n104), .ZN(vscale_core_DW01_add_10n102) );
  INV_X1 vscale_core_DW01_add_10_U400 ( .A(vscale_core_DW01_add_10n143), .ZN(vscale_core_DW01_add_10n289) );
  AND2_X4 vscale_core_DW01_add_10_U401 ( .A1(vscale_core_DW01_add_10n405), .A2(vscale_core_DW01_add_10n277), .ZN(imem_haddr[1]) );
  AOI21_X2 vscale_core_DW01_add_10_U402 ( .B1(vscale_core_DW01_add_10n263), .B2(vscale_core_DW01_add_10n304), .A(vscale_core_DW01_add_10n260), .ZN(vscale_core_DW01_add_10n258) );
  NOR2_X2 vscale_core_DW01_add_10_U403 ( .A1(vscale_core_DW01_add_10n101), .A2(vscale_core_DW01_add_10n135), .ZN(vscale_core_DW01_add_10n4) );
  XNOR2_X2 vscale_core_DW01_add_10_U404 ( .A(vscale_core_DW01_add_10n400), .B(vscale_core_DW01_add_10n409), .ZN(n13174) );
  AND2_X4 vscale_core_DW01_add_10_U405 ( .A1(vscale_core_DW01_add_10n292), .A2(vscale_core_DW01_add_10n165), .ZN(vscale_core_DW01_add_10n400) );
  NAND2_X2 vscale_core_DW01_add_10_U406 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[24]), .ZN(vscale_core_DW01_add_10n106) );
  INV_X1 vscale_core_DW01_add_10_U407 ( .A(vscale_core_DW01_add_10n274), .ZN(vscale_core_DW01_add_10n307) );
  INV_X2 vscale_core_DW01_add_10_U408 ( .A(vscale_core_DW01_add_10n3), .ZN(vscale_core_DW01_add_10n98) );
  NAND2_X2 vscale_core_DW01_add_10_U409 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[25]), .ZN(vscale_core_DW01_add_10n95) );
  INV_X2 vscale_core_DW01_add_10_U410 ( .A(vscale_core_DW01_add_10n204), .ZN(vscale_core_DW01_add_10n206) );
  AOI21_X2 vscale_core_DW01_add_10_U411 ( .B1(vscale_core_DW01_add_10n238), .B2(vscale_core_DW01_add_10n251), .A(vscale_core_DW01_add_10n239), .ZN(vscale_core_DW01_add_10n237) );
  OAI21_X2 vscale_core_DW01_add_10_U412 ( .B1(vscale_core_DW01_add_10n267), .B2(vscale_core_DW01_add_10n271), .A(vscale_core_DW01_add_10n268), .ZN(vscale_core_DW01_add_10n266) );
  AND2_X1 vscale_core_DW01_add_10_U413 ( .A1(pipeline_PCmux_base[11]), .A2(pipeline_PCmux_offset[11]), .ZN(vscale_core_DW01_add_10n401) );
  AOI21_X2 vscale_core_DW01_add_10_U414 ( .B1(vscale_core_DW01_add_10n263), .B2(vscale_core_DW01_add_10n250), .A(vscale_core_DW01_add_10n251), .ZN(vscale_core_DW01_add_10n249) );
  INV_X2 vscale_core_DW01_add_10_U415 ( .A(vscale_core_DW01_add_10n264), .ZN(vscale_core_DW01_add_10n263) );
  OAI21_X2 vscale_core_DW01_add_10_U416 ( .B1(vscale_core_DW01_add_10n234), .B2(vscale_core_DW01_add_10n185), .A(vscale_core_DW01_add_10n186), .ZN(vscale_core_DW01_add_10n184) );
  OAI21_X2 vscale_core_DW01_add_10_U417 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n117), .A(vscale_core_DW01_add_10n118), .ZN(vscale_core_DW01_add_10n116) );
  NOR2_X1 vscale_core_DW01_add_10_U418 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[26]), .ZN(vscale_core_DW01_add_10n402) );
  NOR2_X2 vscale_core_DW01_add_10_U419 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[26]), .ZN(vscale_core_DW01_add_10n87) );
  OAI21_X2 vscale_core_DW01_add_10_U420 ( .B1(vscale_core_DW01_add_10n125), .B2(vscale_core_DW01_add_10n133), .A(vscale_core_DW01_add_10n126), .ZN(vscale_core_DW01_add_10n120) );
  OAI21_X2 vscale_core_DW01_add_10_U421 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n79), .A(vscale_core_DW01_add_10n80), .ZN(vscale_core_DW01_add_10n78) );
  NOR2_X2 vscale_core_DW01_add_10_U422 ( .A1(vscale_core_DW01_add_10n270), .A2(vscale_core_DW01_add_10n267), .ZN(vscale_core_DW01_add_10n265) );
  NAND2_X1 vscale_core_DW01_add_10_U423 ( .A1(pipeline_PCmux_base[16]), .A2(pipeline_PCmux_offset[16]), .ZN(vscale_core_DW01_add_10n174) );
  NOR2_X2 vscale_core_DW01_add_10_U424 ( .A1(pipeline_PCmux_base[13]), .A2(pipeline_PCmux_offset[13]), .ZN(vscale_core_DW01_add_10n200) );
  NOR2_X2 vscale_core_DW01_add_10_U425 ( .A1(vscale_core_DW01_add_10n74), .A2(vscale_core_DW01_add_10n67), .ZN(vscale_core_DW01_add_10n65) );
  AOI21_X2 vscale_core_DW01_add_10_U426 ( .B1(vscale_core_DW01_add_10n263), .B2(vscale_core_DW01_add_10n243), .A(vscale_core_DW01_add_10n244), .ZN(vscale_core_DW01_add_10n242) );
  NOR2_X2 vscale_core_DW01_add_10_U427 ( .A1(pipeline_PCmux_base[11]), .A2(pipeline_PCmux_offset[11]), .ZN(vscale_core_DW01_add_10n218) );
  INV_X1 vscale_core_DW01_add_10_U428 ( .A(vscale_core_DW01_add_10n47), .ZN(vscale_core_DW01_add_10n279) );
  OAI21_X1 vscale_core_DW01_add_10_U429 ( .B1(vscale_core_DW01_add_10n47), .B2(vscale_core_DW01_add_10n57), .A(vscale_core_DW01_add_10n48), .ZN(vscale_core_DW01_add_10n46) );
  OR2_X2 vscale_core_DW01_add_10_U430 ( .A1(vscale_core_DW01_add_10n54), .A2(vscale_core_DW01_add_10n47), .ZN(vscale_core_DW01_add_10n404) );
  NAND2_X1 vscale_core_DW01_add_10_U431 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[30]), .ZN(vscale_core_DW01_add_10n48) );
  NAND2_X2 vscale_core_DW01_add_10_U432 ( .A1(vscale_core_DW01_add_10n411), .A2(pipeline_PCmux_base[28]), .ZN(vscale_core_DW01_add_10n68) );
  NAND2_X2 vscale_core_DW01_add_10_U433 ( .A1(vscale_core_DW01_add_10n4), .A2(vscale_core_DW01_add_10n52), .ZN(vscale_core_DW01_add_10n50) );
  NOR2_X2 vscale_core_DW01_add_10_U434 ( .A1(vscale_core_DW01_add_10n63), .A2(vscale_core_DW01_add_10n54), .ZN(vscale_core_DW01_add_10n52) );
  NOR2_X2 vscale_core_DW01_add_10_U435 ( .A1(pipeline_PCmux_base[16]), .A2(pipeline_PCmux_offset[16]), .ZN(vscale_core_DW01_add_10n173) );
  NOR2_X2 vscale_core_DW01_add_10_U436 ( .A1(pipeline_PCmux_base[15]), .A2(pipeline_PCmux_offset[15]), .ZN(vscale_core_DW01_add_10n180) );
  NAND2_X1 vscale_core_DW01_add_10_U437 ( .A1(vscale_core_DW01_add_10n4), .A2(vscale_core_DW01_add_10n92), .ZN(vscale_core_DW01_add_10n90) );
  NAND2_X1 vscale_core_DW01_add_10_U438 ( .A1(vscale_core_DW01_add_10n4), .A2(vscale_core_DW01_add_10n72), .ZN(vscale_core_DW01_add_10n70) );
  NAND2_X1 vscale_core_DW01_add_10_U439 ( .A1(vscale_core_DW01_add_10n4), .A2(vscale_core_DW01_add_10n61), .ZN(vscale_core_DW01_add_10n59) );
  NAND2_X1 vscale_core_DW01_add_10_U440 ( .A1(vscale_core_DW01_add_10n4), .A2(vscale_core_DW01_add_10n41), .ZN(vscale_core_DW01_add_10n39) );
  NAND2_X1 vscale_core_DW01_add_10_U441 ( .A1(vscale_core_DW01_add_10n4), .A2(vscale_core_DW01_add_10n81), .ZN(vscale_core_DW01_add_10n79) );
  NOR2_X2 vscale_core_DW01_add_10_U442 ( .A1(vscale_core_DW01_add_10n232), .A2(vscale_core_DW01_add_10n229), .ZN(vscale_core_DW01_add_10n223) );
  NOR2_X1 vscale_core_DW01_add_10_U443 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[30]), .ZN(vscale_core_DW01_add_10n47) );
  NAND2_X1 vscale_core_DW01_add_10_U444 ( .A1(vscale_core_DW01_add_10n223), .A2(vscale_core_DW01_add_10n298), .ZN(vscale_core_DW01_add_10n214) );
  INV_X1 vscale_core_DW01_add_10_U445 ( .A(vscale_core_DW01_add_10n223), .ZN(vscale_core_DW01_add_10n221) );
  NAND2_X2 vscale_core_DW01_add_10_U446 ( .A1(vscale_core_DW01_add_10n297), .A2(vscale_core_DW01_add_10n212), .ZN(vscale_core_DW01_add_10n24) );
  NAND2_X2 vscale_core_DW01_add_10_U447 ( .A1(vscale_core_DW01_add_10n293), .A2(vscale_core_DW01_add_10n174), .ZN(vscale_core_DW01_add_10n20) );
  NAND2_X2 vscale_core_DW01_add_10_U448 ( .A1(vscale_core_DW01_add_10n299), .A2(vscale_core_DW01_add_10n230), .ZN(vscale_core_DW01_add_10n26) );
  NAND2_X2 vscale_core_DW01_add_10_U449 ( .A1(vscale_core_DW01_add_10n296), .A2(vscale_core_DW01_add_10n201), .ZN(vscale_core_DW01_add_10n23) );
  NAND2_X2 vscale_core_DW01_add_10_U450 ( .A1(vscale_core_DW01_add_10n294), .A2(vscale_core_DW01_add_10n183), .ZN(vscale_core_DW01_add_10n21) );
  NAND2_X2 vscale_core_DW01_add_10_U451 ( .A1(vscale_core_DW01_add_10n301), .A2(vscale_core_DW01_add_10n241), .ZN(vscale_core_DW01_add_10n28) );
  NOR2_X1 vscale_core_DW01_add_10_U452 ( .A1(pipeline_PCmux_base[9]), .A2(pipeline_PCmux_offset[9]), .ZN(vscale_core_DW01_add_10n232) );
  INV_X1 vscale_core_DW01_add_10_U453 ( .A(vscale_core_DW01_add_10n224), .ZN(vscale_core_DW01_add_10n222) );
  NOR2_X1 vscale_core_DW01_add_10_U454 ( .A1(vscale_core_DW01_add_10n121), .A2(vscale_core_DW01_add_10n112), .ZN(vscale_core_DW01_add_10n110) );
  INV_X1 vscale_core_DW01_add_10_U455 ( .A(vscale_core_DW01_add_10n267), .ZN(vscale_core_DW01_add_10n305) );
  XOR2_X2 vscale_core_DW01_add_10_U456 ( .A(vscale_core_DW01_add_10n403), .B(vscale_core_DW01_add_10n272), .Z(imem_haddr[3]) );
  NAND2_X1 vscale_core_DW01_add_10_U457 ( .A1(vscale_core_DW01_add_10n306), .A2(vscale_core_DW01_add_10n271), .ZN(vscale_core_DW01_add_10n403) );
  AOI21_X1 vscale_core_DW01_add_10_U458 ( .B1(vscale_core_DW01_add_10n206), .B2(vscale_core_DW01_add_10n178), .A(vscale_core_DW01_add_10n179), .ZN(vscale_core_DW01_add_10n177) );
  AOI21_X1 vscale_core_DW01_add_10_U459 ( .B1(vscale_core_DW01_add_10n206), .B2(vscale_core_DW01_add_10n296), .A(vscale_core_DW01_add_10n199), .ZN(vscale_core_DW01_add_10n197) );
  OAI21_X1 vscale_core_DW01_add_10_U460 ( .B1(vscale_core_DW01_add_10n253), .B2(vscale_core_DW01_add_10n245), .A(vscale_core_DW01_add_10n248), .ZN(vscale_core_DW01_add_10n244) );
  NOR2_X1 vscale_core_DW01_add_10_U461 ( .A1(vscale_core_DW01_add_10n252), .A2(vscale_core_DW01_add_10n245), .ZN(vscale_core_DW01_add_10n243) );
  INV_X1 vscale_core_DW01_add_10_U462 ( .A(vscale_core_DW01_add_10n82), .ZN(vscale_core_DW01_add_10n84) );
  INV_X1 vscale_core_DW01_add_10_U463 ( .A(vscale_core_DW01_add_10n151), .ZN(vscale_core_DW01_add_10n149) );
  NAND2_X1 vscale_core_DW01_add_10_U464 ( .A1(vscale_core_DW01_add_10n300), .A2(vscale_core_DW01_add_10n233), .ZN(vscale_core_DW01_add_10n27) );
  NOR2_X1 vscale_core_DW01_add_10_U465 ( .A1(vscale_core_DW01_add_10n83), .A2(vscale_core_DW01_add_10n74), .ZN(vscale_core_DW01_add_10n72) );
  NAND2_X1 vscale_core_DW01_add_10_U466 ( .A1(vscale_core_DW01_add_10n302), .A2(vscale_core_DW01_add_10n248), .ZN(vscale_core_DW01_add_10n29) );
  INV_X4 vscale_core_DW01_add_10_U467 ( .A(n6781), .ZN(vscale_core_DW01_add_10n412) );
  OAI21_X1 vscale_core_DW01_add_10_U468 ( .B1(vscale_core_DW01_add_10n234), .B2(vscale_core_DW01_add_10n203), .A(vscale_core_DW01_add_10n204), .ZN(vscale_core_DW01_add_10n202) );
  AOI21_X1 vscale_core_DW01_add_10_U469 ( .B1(vscale_core_DW01_add_10n138), .B2(vscale_core_DW01_add_10n119), .A(vscale_core_DW01_add_10n120), .ZN(vscale_core_DW01_add_10n118) );
  AOI21_X1 vscale_core_DW01_add_10_U470 ( .B1(vscale_core_DW01_add_10n206), .B2(vscale_core_DW01_add_10n187), .A(vscale_core_DW01_add_10n188), .ZN(vscale_core_DW01_add_10n186) );
  OAI21_X1 vscale_core_DW01_add_10_U471 ( .B1(vscale_core_DW01_add_10n234), .B2(vscale_core_DW01_add_10n221), .A(vscale_core_DW01_add_10n222), .ZN(vscale_core_DW01_add_10n220) );
  NOR2_X2 vscale_core_DW01_add_10_U472 ( .A1(vscale_core_DW01_add_10n63), .A2(vscale_core_DW01_add_10n404), .ZN(vscale_core_DW01_add_10n41) );
  OAI21_X1 vscale_core_DW01_add_10_U473 ( .B1(vscale_core_DW01_add_10n272), .B2(vscale_core_DW01_add_10n270), .A(vscale_core_DW01_add_10n271), .ZN(vscale_core_DW01_add_10n269) );
  OAI21_X2 vscale_core_DW01_add_10_U474 ( .B1(vscale_core_DW01_add_10n105), .B2(vscale_core_DW01_add_10n115), .A(vscale_core_DW01_add_10n106), .ZN(vscale_core_DW01_add_10n104) );
  OAI21_X2 vscale_core_DW01_add_10_U475 ( .B1(vscale_core_DW01_add_10n143), .B2(vscale_core_DW01_add_10n151), .A(vscale_core_DW01_add_10n144), .ZN(vscale_core_DW01_add_10n142) );
  NOR2_X2 vscale_core_DW01_add_10_U476 ( .A1(vscale_core_DW01_add_10n245), .A2(vscale_core_DW01_add_10n240), .ZN(vscale_core_DW01_add_10n238) );
  OAI21_X1 vscale_core_DW01_add_10_U477 ( .B1(vscale_core_DW01_add_10n84), .B2(vscale_core_DW01_add_10n74), .A(vscale_core_DW01_add_10n77), .ZN(vscale_core_DW01_add_10n73) );
  OAI21_X2 vscale_core_DW01_add_10_U478 ( .B1(vscale_core_DW01_add_10n240), .B2(vscale_core_DW01_add_10n248), .A(vscale_core_DW01_add_10n241), .ZN(vscale_core_DW01_add_10n239) );
  OAI21_X1 vscale_core_DW01_add_10_U479 ( .B1(vscale_core_DW01_add_10n122), .B2(vscale_core_DW01_add_10n112), .A(vscale_core_DW01_add_10n115), .ZN(vscale_core_DW01_add_10n111) );
  OAI21_X1 vscale_core_DW01_add_10_U480 ( .B1(vscale_core_DW01_add_10n190), .B2(vscale_core_DW01_add_10n180), .A(vscale_core_DW01_add_10n183), .ZN(vscale_core_DW01_add_10n179) );
  OAI21_X1 vscale_core_DW01_add_10_U481 ( .B1(vscale_core_DW01_add_10n234), .B2(vscale_core_DW01_add_10n232), .A(vscale_core_DW01_add_10n233), .ZN(vscale_core_DW01_add_10n231) );
  AOI21_X1 vscale_core_DW01_add_10_U482 ( .B1(vscale_core_DW01_add_10n156), .B2(vscale_core_DW01_add_10n290), .A(vscale_core_DW01_add_10n149), .ZN(vscale_core_DW01_add_10n147) );
  OAI21_X1 vscale_core_DW01_add_10_U483 ( .B1(vscale_core_DW01_add_10n234), .B2(vscale_core_DW01_add_10n214), .A(vscale_core_DW01_add_10n215), .ZN(vscale_core_DW01_add_10n213) );
  OAI21_X1 vscale_core_DW01_add_10_U484 ( .B1(vscale_core_DW01_add_10n234), .B2(vscale_core_DW01_add_10n176), .A(vscale_core_DW01_add_10n177), .ZN(vscale_core_DW01_add_10n175) );
  NOR2_X1 vscale_core_DW01_add_10_U485 ( .A1(vscale_core_DW01_add_10n189), .A2(vscale_core_DW01_add_10n180), .ZN(vscale_core_DW01_add_10n178) );
  OAI21_X1 vscale_core_DW01_add_10_U486 ( .B1(vscale_core_DW01_add_10n234), .B2(vscale_core_DW01_add_10n196), .A(vscale_core_DW01_add_10n197), .ZN(vscale_core_DW01_add_10n195) );
  NOR2_X2 vscale_core_DW01_add_10_U487 ( .A1(vscale_core_DW01_add_10n164), .A2(vscale_core_DW01_add_10n161), .ZN(vscale_core_DW01_add_10n155) );
  OAI21_X2 vscale_core_DW01_add_10_U488 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n50), .A(vscale_core_DW01_add_10n51), .ZN(vscale_core_DW01_add_10n49) );
  OAI21_X2 vscale_core_DW01_add_10_U489 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n39), .A(vscale_core_DW01_add_10n40), .ZN(vscale_core_DW01_add_10n38) );
  INV_X4 vscale_core_DW01_add_10_U490 ( .A(vscale_core_DW01_add_10n412), .ZN(vscale_core_DW01_add_10n410) );
  INV_X4 vscale_core_DW01_add_10_U491 ( .A(vscale_core_DW01_add_10n412), .ZN(vscale_core_DW01_add_10n411) );
  OR2_X1 vscale_core_DW01_add_10_U492 ( .A1(pipeline_PCmux_base[1]), .A2(pipeline_PCmux_offset[1]), .ZN(vscale_core_DW01_add_10n405) );
  NOR2_X2 vscale_core_DW01_add_10_U493 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[23]), .ZN(vscale_core_DW01_add_10n112) );
  NOR2_X2 vscale_core_DW01_add_10_U494 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[27]), .ZN(vscale_core_DW01_add_10n74) );
  NOR2_X2 vscale_core_DW01_add_10_U495 ( .A1(pipeline_PCmux_base[7]), .A2(pipeline_PCmux_offset[7]), .ZN(vscale_core_DW01_add_10n245) );
  NOR2_X2 vscale_core_DW01_add_10_U496 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[29]), .ZN(vscale_core_DW01_add_10n54) );
  NOR2_X2 vscale_core_DW01_add_10_U497 ( .A1(pipeline_PCmux_base[3]), .A2(pipeline_PCmux_offset[3]), .ZN(vscale_core_DW01_add_10n270) );
  NAND2_X2 vscale_core_DW01_add_10_U498 ( .A1(pipeline_PCmux_base[19]), .A2(pipeline_PCmux_offset[19]), .ZN(vscale_core_DW01_add_10n151) );
  NOR2_X1 vscale_core_DW01_add_10_U499 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[25]), .ZN(vscale_core_DW01_add_10n94) );
  NAND2_X2 vscale_core_DW01_add_10_U500 ( .A1(pipeline_PCmux_base[11]), .A2(pipeline_PCmux_offset[11]), .ZN(vscale_core_DW01_add_10n219) );
  OR2_X1 vscale_core_DW01_add_10_U501 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[31]), .ZN(vscale_core_DW01_add_10n406) );
  BUF_X4 vscale_core_DW01_add_10_U502 ( .A(pipeline_PCmux_base[0]), .Z(imem_haddr[0]) );
  NOR2_X2 vscale_core_DW01_add_10_U503 ( .A1(vscale_core_DW01_add_10n94), .A2(vscale_core_DW01_add_10n402), .ZN(vscale_core_DW01_add_10n81) );
  INV_X1 vscale_core_DW01_add_10_U504 ( .A(vscale_core_DW01_add_10n402), .ZN(vscale_core_DW01_add_10n283) );
  AOI21_X2 vscale_core_DW01_add_10_U505 ( .B1(vscale_core_DW01_add_10n224), .B2(vscale_core_DW01_add_10n298), .A(vscale_core_DW01_add_10n401), .ZN(vscale_core_DW01_add_10n215) );
  NOR2_X2 vscale_core_DW01_add_10_U506 ( .A1(vscale_core_DW01_add_10n143), .A2(vscale_core_DW01_add_10n150), .ZN(vscale_core_DW01_add_10n141) );
  OAI21_X2 vscale_core_DW01_add_10_U507 ( .B1(vscale_core_DW01_add_10n67), .B2(vscale_core_DW01_add_10n77), .A(vscale_core_DW01_add_10n68), .ZN(vscale_core_DW01_add_10n66) );
  OAI21_X2 vscale_core_DW01_add_10_U508 ( .B1(vscale_core_DW01_add_10n87), .B2(vscale_core_DW01_add_10n95), .A(vscale_core_DW01_add_10n88), .ZN(vscale_core_DW01_add_10n82) );
  OAI21_X2 vscale_core_DW01_add_10_U509 ( .B1(vscale_core_DW01_add_10n173), .B2(vscale_core_DW01_add_10n183), .A(vscale_core_DW01_add_10n174), .ZN(vscale_core_DW01_add_10n172) );
  INV_X1 vscale_core_DW01_add_10_U510 ( .A(vscale_core_DW01_add_10n173), .ZN(vscale_core_DW01_add_10n293) );
  OAI21_X2 vscale_core_DW01_add_10_U511 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n70), .A(vscale_core_DW01_add_10n71), .ZN(vscale_core_DW01_add_10n69) );
  OAI21_X2 vscale_core_DW01_add_10_U512 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n59), .A(vscale_core_DW01_add_10n60), .ZN(vscale_core_DW01_add_10n58) );
  OAI21_X2 vscale_core_DW01_add_10_U513 ( .B1(vscale_core_DW01_add_10n409), .B2(vscale_core_DW01_add_10n90), .A(vscale_core_DW01_add_10n91), .ZN(vscale_core_DW01_add_10n89) );
  INV_X1 vscale_core_DW01_add_10_U514 ( .A(vscale_core_DW01_add_10n125), .ZN(vscale_core_DW01_add_10n287) );
  NAND2_X1 vscale_core_DW01_add_10_U515 ( .A1(vscale_core_DW01_add_10n298), .A2(vscale_core_DW01_add_10n219), .ZN(vscale_core_DW01_add_10n25) );
  NOR2_X2 vscale_core_DW01_add_10_U516 ( .A1(vscale_core_DW01_add_10n218), .A2(vscale_core_DW01_add_10n211), .ZN(vscale_core_DW01_add_10n209) );
  NOR2_X2 vscale_core_DW01_add_10_U517 ( .A1(pipeline_PCmux_base[19]), .A2(pipeline_PCmux_offset[19]), .ZN(vscale_core_DW01_add_10n150) );
  XOR2_X2 vscale_core_DW01_add_10_U518 ( .A(vscale_core_DW01_add_10n27), .B(vscale_core_DW01_add_10n234), .Z(n13182) );
  OAI21_X2 vscale_core_DW01_add_10_U519 ( .B1(vscale_core_DW01_add_10n64), .B2(vscale_core_DW01_add_10n54), .A(vscale_core_DW01_add_10n57), .ZN(vscale_core_DW01_add_10n53) );
  OAI21_X2 vscale_core_DW01_add_10_U520 ( .B1(vscale_core_DW01_add_10n64), .B2(vscale_core_DW01_add_10n404), .A(vscale_core_DW01_add_10n44), .ZN(vscale_core_DW01_add_10n42) );
  INV_X1 vscale_core_DW01_add_10_U521 ( .A(vscale_core_DW01_add_10n64), .ZN(vscale_core_DW01_add_10n62) );
  NOR2_X2 vscale_core_DW01_add_10_U522 ( .A1(vscale_core_DW01_add_10n410), .A2(pipeline_PCmux_base[21]), .ZN(vscale_core_DW01_add_10n132) );
  AOI21_X2 vscale_core_DW01_add_10_U523 ( .B1(vscale_core_DW01_add_10n3), .B2(vscale_core_DW01_add_10n81), .A(vscale_core_DW01_add_10n82), .ZN(vscale_core_DW01_add_10n80) );
  AOI21_X2 vscale_core_DW01_add_10_U524 ( .B1(vscale_core_DW01_add_10n3), .B2(vscale_core_DW01_add_10n92), .A(vscale_core_DW01_add_10n93), .ZN(vscale_core_DW01_add_10n91) );
  AOI21_X2 vscale_core_DW01_add_10_U525 ( .B1(vscale_core_DW01_add_10n3), .B2(vscale_core_DW01_add_10n72), .A(vscale_core_DW01_add_10n73), .ZN(vscale_core_DW01_add_10n71) );
  AOI21_X2 vscale_core_DW01_add_10_U526 ( .B1(vscale_core_DW01_add_10n3), .B2(vscale_core_DW01_add_10n61), .A(vscale_core_DW01_add_10n62), .ZN(vscale_core_DW01_add_10n60) );
  OAI21_X2 vscale_core_DW01_add_10_U527 ( .B1(vscale_core_DW01_add_10n204), .B2(vscale_core_DW01_add_10n169), .A(vscale_core_DW01_add_10n170), .ZN(vscale_core_DW01_add_10n168) );
  INV_X4 vscale_core_DW01_add_10_U528 ( .A(vscale_core_DW01_add_10n4), .ZN(vscale_core_DW01_add_10n97) );
  INV_X4 vscale_core_DW01_add_10_U529 ( .A(vscale_core_DW01_add_10n95), .ZN(vscale_core_DW01_add_10n93) );
  INV_X4 vscale_core_DW01_add_10_U530 ( .A(vscale_core_DW01_add_10n81), .ZN(vscale_core_DW01_add_10n83) );
  INV_X4 vscale_core_DW01_add_10_U531 ( .A(vscale_core_DW01_add_10n63), .ZN(vscale_core_DW01_add_10n61) );
  INV_X4 vscale_core_DW01_add_10_U532 ( .A(vscale_core_DW01_add_10n46), .ZN(vscale_core_DW01_add_10n44) );
  INV_X4 vscale_core_DW01_add_10_U533 ( .A(vscale_core_DW01_add_10n270), .ZN(vscale_core_DW01_add_10n306) );
  INV_X4 vscale_core_DW01_add_10_U534 ( .A(vscale_core_DW01_add_10n245), .ZN(vscale_core_DW01_add_10n302) );
  INV_X4 vscale_core_DW01_add_10_U535 ( .A(vscale_core_DW01_add_10n240), .ZN(vscale_core_DW01_add_10n301) );
  INV_X4 vscale_core_DW01_add_10_U536 ( .A(vscale_core_DW01_add_10n232), .ZN(vscale_core_DW01_add_10n300) );
  INV_X4 vscale_core_DW01_add_10_U537 ( .A(vscale_core_DW01_add_10n229), .ZN(vscale_core_DW01_add_10n299) );
  INV_X4 vscale_core_DW01_add_10_U538 ( .A(vscale_core_DW01_add_10n211), .ZN(vscale_core_DW01_add_10n297) );
  INV_X4 vscale_core_DW01_add_10_U539 ( .A(vscale_core_DW01_add_10n193), .ZN(vscale_core_DW01_add_10n295) );
  INV_X4 vscale_core_DW01_add_10_U540 ( .A(vscale_core_DW01_add_10n180), .ZN(vscale_core_DW01_add_10n294) );
  INV_X4 vscale_core_DW01_add_10_U541 ( .A(vscale_core_DW01_add_10n164), .ZN(vscale_core_DW01_add_10n292) );
  INV_X4 vscale_core_DW01_add_10_U542 ( .A(vscale_core_DW01_add_10n161), .ZN(vscale_core_DW01_add_10n291) );
  INV_X4 vscale_core_DW01_add_10_U543 ( .A(vscale_core_DW01_add_10n112), .ZN(vscale_core_DW01_add_10n286) );
  INV_X4 vscale_core_DW01_add_10_U544 ( .A(vscale_core_DW01_add_10n105), .ZN(vscale_core_DW01_add_10n285) );
  INV_X4 vscale_core_DW01_add_10_U545 ( .A(vscale_core_DW01_add_10n94), .ZN(vscale_core_DW01_add_10n92) );
  INV_X4 vscale_core_DW01_add_10_U546 ( .A(vscale_core_DW01_add_10n74), .ZN(vscale_core_DW01_add_10n282) );
  INV_X4 vscale_core_DW01_add_10_U547 ( .A(vscale_core_DW01_add_10n67), .ZN(vscale_core_DW01_add_10n281) );
  INV_X4 vscale_core_DW01_add_10_U548 ( .A(vscale_core_DW01_add_10n54), .ZN(vscale_core_DW01_add_10n280) );
  INV_X4 vscale_core_DW01_add_10_U549 ( .A(vscale_core_DW01_add_10n262), .ZN(vscale_core_DW01_add_10n260) );
  INV_X4 vscale_core_DW01_add_10_U550 ( .A(vscale_core_DW01_add_10n261), .ZN(vscale_core_DW01_add_10n304) );
  INV_X4 vscale_core_DW01_add_10_U551 ( .A(vscale_core_DW01_add_10n251), .ZN(vscale_core_DW01_add_10n253) );
  INV_X4 vscale_core_DW01_add_10_U552 ( .A(vscale_core_DW01_add_10n250), .ZN(vscale_core_DW01_add_10n252) );
  INV_X4 vscale_core_DW01_add_10_U553 ( .A(vscale_core_DW01_add_10n235), .ZN(vscale_core_DW01_add_10n234) );
  INV_X4 vscale_core_DW01_add_10_U554 ( .A(vscale_core_DW01_add_10n218), .ZN(vscale_core_DW01_add_10n298) );
  INV_X4 vscale_core_DW01_add_10_U555 ( .A(vscale_core_DW01_add_10n203), .ZN(vscale_core_DW01_add_10n205) );
  INV_X4 vscale_core_DW01_add_10_U556 ( .A(vscale_core_DW01_add_10n201), .ZN(vscale_core_DW01_add_10n199) );
  INV_X4 vscale_core_DW01_add_10_U557 ( .A(vscale_core_DW01_add_10n200), .ZN(vscale_core_DW01_add_10n296) );
  INV_X4 vscale_core_DW01_add_10_U558 ( .A(vscale_core_DW01_add_10n188), .ZN(vscale_core_DW01_add_10n190) );
  INV_X4 vscale_core_DW01_add_10_U559 ( .A(vscale_core_DW01_add_10n187), .ZN(vscale_core_DW01_add_10n189) );
  INV_X4 vscale_core_DW01_add_10_U560 ( .A(vscale_core_DW01_add_10n156), .ZN(vscale_core_DW01_add_10n154) );
  INV_X4 vscale_core_DW01_add_10_U561 ( .A(vscale_core_DW01_add_10n155), .ZN(vscale_core_DW01_add_10n153) );
  INV_X4 vscale_core_DW01_add_10_U562 ( .A(vscale_core_DW01_add_10n150), .ZN(vscale_core_DW01_add_10n290) );
  INV_X4 vscale_core_DW01_add_10_U563 ( .A(vscale_core_DW01_add_10n136), .ZN(vscale_core_DW01_add_10n138) );
  INV_X4 vscale_core_DW01_add_10_U564 ( .A(vscale_core_DW01_add_10n135), .ZN(vscale_core_DW01_add_10n137) );
  INV_X4 vscale_core_DW01_add_10_U565 ( .A(vscale_core_DW01_add_10n133), .ZN(vscale_core_DW01_add_10n131) );
  INV_X4 vscale_core_DW01_add_10_U566 ( .A(vscale_core_DW01_add_10n132), .ZN(vscale_core_DW01_add_10n288) );
  INV_X4 vscale_core_DW01_add_10_U567 ( .A(vscale_core_DW01_add_10n120), .ZN(vscale_core_DW01_add_10n122) );
  INV_X4 vscale_core_DW01_add_10_U568 ( .A(vscale_core_DW01_add_10n119), .ZN(vscale_core_DW01_add_10n121) );
;


  DFF_X1 pipeline_md_b_reg_5_ ( .D(n5775), .CK(clk), .Q(pipeline_md_b[5]), 
        .QN(n6919) );
  DFF_X1 pipeline_md_b_reg_4_ ( .D(n5776), .CK(clk), .Q(pipeline_md_b[4]), 
        .QN(n6718) );
  DFF_X1 pipeline_md_b_reg_3_ ( .D(n5777), .CK(clk), .Q(pipeline_md_b[3]), 
        .QN(n6760) );
  DFF_X1 pipeline_md_b_reg_2_ ( .D(n5778), .CK(clk), .Q(pipeline_md_b[2]), 
        .QN(n6920) );
  DFF_X1 pipeline_md_b_reg_1_ ( .D(n5779), .CK(clk), .Q(pipeline_md_b[1]), 
        .QN(n6759) );
  DFF_X1 pipeline_md_b_reg_0_ ( .D(n5780), .CK(clk), .Q(pipeline_md_b[0]), 
        .QN(n6921) );
  DFF_X2 pipeline_md_a_reg_31_ ( .D(n5684), .CK(clk), .Q(pipeline_md_a[31]), 
        .QN(n13057) );
  DFF_X2 pipeline_md_a_reg_30_ ( .D(n5683), .CK(clk), .Q(pipeline_md_a[30]), 
        .QN(n13058) );
  DFF_X2 pipeline_md_a_reg_58_ ( .D(n5711), .CK(clk), .Q(pipeline_md_a[58]), 
        .QN(n1145) );
  DFF_X2 pipeline_md_a_reg_59_ ( .D(n5712), .CK(clk), .Q(pipeline_md_a[59]), 
        .QN(n1146) );
  DFF_X2 pipeline_md_a_reg_60_ ( .D(n5713), .CK(clk), .Q(pipeline_md_a[60]), 
        .QN(n1147) );
  DFF_X2 pipeline_md_a_reg_61_ ( .D(n5714), .CK(clk), .Q(pipeline_md_a[61]), 
        .QN(n1148) );
  DFF_X1 pipeline_ctrl_replay_IF_reg ( .D(pipeline_ctrl_N66), .CK(clk), .Q(
        pipeline_ctrl_replay_IF), .QN(n6922) );
  DFF_X1 pipeline_inst_DX_reg_1_ ( .D(n6256), .CK(clk), .Q(pipeline_inst_DX[1]) );
  DFF_X1 pipeline_inst_DX_reg_0_ ( .D(n6294), .CK(clk), .Q(pipeline_inst_DX[0]) );
  DFF_X1 pipeline_md_counter_reg_1_ ( .D(n6250), .CK(clk), .Q(pipeline_md_N22), 
        .QN(n6747) );
  DFF_X1 pipeline_md_state_reg_0_ ( .D(pipeline_md_N161), .CK(clk), .Q(
        pipeline_md_state[0]), .QN(n6810) );
  DFF_X2 pipeline_csr_mtvec_reg_31_ ( .D(n6177), .CK(clk), .Q(n10282), .QN(
        n1222) );
  DFF_X2 pipeline_md_result_reg_58_ ( .D(n5595), .CK(clk), .Q(
        pipeline_md_result[58]), .QN(n950) );
  DFF_X2 pipeline_md_result_reg_59_ ( .D(n5594), .CK(clk), .Q(
        pipeline_md_result[59]), .QN(n952) );
  DFF_X2 pipeline_md_result_reg_60_ ( .D(n5593), .CK(clk), .Q(
        pipeline_md_result[60]), .QN(n954) );
  DFF_X1 pipeline_csr_cycle_full_reg_7_ ( .D(pipeline_csr_N1895), .CK(clk), 
        .Q(pipeline_csr_cycle_full[7]) );
  DFF_X1 pipeline_csr_cycle_full_reg_0_ ( .D(pipeline_csr_N1888), .CK(clk), 
        .Q(pipeline_csr_cycle_full[0]) );
  DFF_X1 pipeline_csr_cycle_full_reg_3_ ( .D(pipeline_csr_N1891), .CK(clk), 
        .Q(pipeline_csr_cycle_full[3]) );
  DFF_X1 pipeline_csr_cycle_full_reg_28_ ( .D(pipeline_csr_N1916), .CK(clk), 
        .Q(pipeline_csr_cycle_full[28]), .QN(n6752) );
  DFF_X1 pipeline_csr_cycle_full_reg_31_ ( .D(pipeline_csr_N1919), .CK(clk), 
        .Q(pipeline_csr_cycle_full[31]), .QN(n6838) );
  DFF_X1 pipeline_csr_cycle_full_reg_32_ ( .D(pipeline_csr_N1920), .CK(clk), 
        .Q(pipeline_csr_cycle_full[32]), .QN(n6829) );
  DFF_X1 pipeline_csr_cycle_full_reg_35_ ( .D(pipeline_csr_N1923), .CK(clk), 
        .Q(pipeline_csr_cycle_full[35]) );
  DFF_X1 pipeline_csr_cycle_full_reg_39_ ( .D(pipeline_csr_N1927), .CK(clk), 
        .Q(pipeline_csr_cycle_full[39]), .QN(n6845) );
  DFF_X1 pipeline_csr_cycle_full_reg_60_ ( .D(pipeline_csr_N1948), .CK(clk), 
        .Q(pipeline_csr_cycle_full[60]), .QN(n6869) );
  DFF_X1 pipeline_csr_cycle_full_reg_62_ ( .D(pipeline_csr_N1950), .CK(clk), 
        .Q(pipeline_csr_cycle_full[62]), .QN(n6866) );
  DFF_X1 pipeline_csr_time_full_reg_30_ ( .D(pipeline_csr_N1982), .CK(clk), 
        .Q(pipeline_csr_time_full[30]), .QN(n6830) );
  DFF_X1 pipeline_csr_time_full_reg_0_ ( .D(pipeline_csr_N1952), .CK(clk), .Q(
        pipeline_csr_time_full[0]) );
  DFF_X1 pipeline_csr_time_full_reg_3_ ( .D(pipeline_csr_N1955), .CK(clk), .Q(
        pipeline_csr_time_full[3]), .QN(n6839) );
  DFF_X1 pipeline_csr_time_full_reg_7_ ( .D(pipeline_csr_N1959), .CK(clk), .Q(
        pipeline_csr_time_full[7]), .QN(n6842) );
  DFF_X1 pipeline_csr_time_full_reg_28_ ( .D(pipeline_csr_N1980), .CK(clk), 
        .Q(pipeline_csr_time_full[28]), .QN(n6831) );
  DFF_X1 pipeline_csr_time_full_reg_31_ ( .D(pipeline_csr_N1983), .CK(clk), 
        .Q(pipeline_csr_time_full[31]), .QN(n6897) );
  DFF_X1 pipeline_csr_time_full_reg_32_ ( .D(pipeline_csr_N1984), .CK(clk), 
        .Q(pipeline_csr_time_full[32]) );
  DFF_X1 pipeline_csr_time_full_reg_35_ ( .D(pipeline_csr_N1987), .CK(clk), 
        .Q(pipeline_csr_time_full[35]), .QN(n6837) );
  DFF_X1 pipeline_csr_time_full_reg_39_ ( .D(pipeline_csr_N1991), .CK(clk), 
        .Q(pipeline_csr_time_full[39]) );
  DFF_X1 pipeline_csr_time_full_reg_60_ ( .D(pipeline_csr_N2012), .CK(clk), 
        .Q(pipeline_csr_time_full[60]) );
  DFF_X1 pipeline_csr_time_full_reg_61_ ( .D(pipeline_csr_N2013), .CK(clk), 
        .Q(pipeline_csr_time_full[61]), .QN(n6868) );
  DFF_X1 pipeline_csr_mtime_full_reg_29_ ( .D(pipeline_csr_N2130), .CK(clk), 
        .Q(pipeline_csr_mtime_full[29]) );
  DFF_X1 pipeline_csr_mtime_full_reg_0_ ( .D(pipeline_csr_N2101), .CK(clk), 
        .Q(pipeline_csr_mtime_full[0]), .QN(n6823) );
  DFF_X1 pipeline_csr_mtime_full_reg_3_ ( .D(pipeline_csr_N2104), .CK(clk), 
        .Q(pipeline_csr_mtime_full[3]) );
  DFF_X1 pipeline_csr_mtime_full_reg_7_ ( .D(pipeline_csr_N2108), .CK(clk), 
        .Q(pipeline_csr_mtime_full[7]), .QN(n6861) );
  DFF_X1 pipeline_csr_mtime_full_reg_28_ ( .D(pipeline_csr_N2129), .CK(clk), 
        .Q(pipeline_csr_mtime_full[28]) );
  DFF_X1 pipeline_csr_mtime_full_reg_30_ ( .D(pipeline_csr_N2131), .CK(clk), 
        .Q(pipeline_csr_mtime_full[30]) );
  DFF_X1 pipeline_csr_mtime_full_reg_31_ ( .D(pipeline_csr_N2132), .CK(clk), 
        .Q(pipeline_csr_mtime_full[31]), .QN(n6828) );
  DFF_X1 pipeline_csr_mtime_full_reg_32_ ( .D(pipeline_csr_N2133), .CK(clk), 
        .Q(pipeline_csr_mtime_full[32]), .QN(n6834) );
  DFF_X1 pipeline_csr_mtime_full_reg_35_ ( .D(pipeline_csr_N2136), .CK(clk), 
        .Q(pipeline_csr_mtime_full[35]) );
  DFF_X1 pipeline_csr_mtime_full_reg_39_ ( .D(pipeline_csr_N2140), .CK(clk), 
        .Q(pipeline_csr_mtime_full[39]), .QN(n6841) );
  DFF_X1 pipeline_csr_mtime_full_reg_59_ ( .D(pipeline_csr_N2160), .CK(clk), 
        .Q(pipeline_csr_mtime_full[59]), .QN(n6870) );
  DFF_X1 pipeline_csr_mtime_full_reg_27_ ( .D(pipeline_csr_N2128), .CK(clk), 
        .Q(pipeline_csr_mtime_full[27]), .QN(n6862) );
  DFF_X1 pipeline_csr_time_full_reg_59_ ( .D(pipeline_csr_N2011), .CK(clk), 
        .Q(pipeline_csr_time_full[59]), .QN(n6871) );
  DFF_X1 pipeline_csr_time_full_reg_27_ ( .D(pipeline_csr_N1979), .CK(clk), 
        .Q(pipeline_csr_time_full[27]), .QN(n6898) );
  DFF_X1 pipeline_csr_cycle_full_reg_59_ ( .D(pipeline_csr_N1947), .CK(clk), 
        .Q(pipeline_csr_cycle_full[59]) );
  DFF_X1 pipeline_csr_cycle_full_reg_27_ ( .D(pipeline_csr_N1915), .CK(clk), 
        .Q(pipeline_csr_cycle_full[27]) );
  DFF_X1 pipeline_csr_mtime_full_reg_58_ ( .D(pipeline_csr_N2159), .CK(clk), 
        .Q(pipeline_csr_mtime_full[58]), .QN(n6872) );
  DFF_X1 pipeline_csr_mtime_full_reg_26_ ( .D(pipeline_csr_N2127), .CK(clk), 
        .Q(pipeline_csr_mtime_full[26]) );
  DFF_X1 pipeline_csr_time_full_reg_58_ ( .D(pipeline_csr_N2010), .CK(clk), 
        .Q(pipeline_csr_time_full[58]), .QN(n6873) );
  DFF_X1 pipeline_csr_time_full_reg_26_ ( .D(pipeline_csr_N1978), .CK(clk), 
        .Q(pipeline_csr_time_full[26]), .QN(n6832) );
  DFF_X1 pipeline_csr_cycle_full_reg_58_ ( .D(pipeline_csr_N1946), .CK(clk), 
        .Q(pipeline_csr_cycle_full[58]) );
  DFF_X1 pipeline_csr_cycle_full_reg_26_ ( .D(pipeline_csr_N1914), .CK(clk), 
        .Q(pipeline_csr_cycle_full[26]) );
  DFF_X1 pipeline_csr_mtime_full_reg_57_ ( .D(pipeline_csr_N2158), .CK(clk), 
        .Q(pipeline_csr_mtime_full[57]), .QN(n6874) );
  DFF_X1 pipeline_csr_mtime_full_reg_25_ ( .D(pipeline_csr_N2126), .CK(clk), 
        .Q(pipeline_csr_mtime_full[25]) );
  DFF_X1 pipeline_csr_time_full_reg_57_ ( .D(pipeline_csr_N2009), .CK(clk), 
        .Q(pipeline_csr_time_full[57]), .QN(n6875) );
  DFF_X1 pipeline_csr_time_full_reg_25_ ( .D(pipeline_csr_N1977), .CK(clk), 
        .Q(pipeline_csr_time_full[25]), .QN(n6899) );
  DFF_X1 pipeline_csr_cycle_full_reg_57_ ( .D(pipeline_csr_N1945), .CK(clk), 
        .Q(pipeline_csr_cycle_full[57]) );
  DFF_X1 pipeline_csr_cycle_full_reg_25_ ( .D(pipeline_csr_N1913), .CK(clk), 
        .Q(pipeline_csr_cycle_full[25]) );
  DFF_X1 pipeline_csr_mtime_full_reg_56_ ( .D(pipeline_csr_N2157), .CK(clk), 
        .Q(pipeline_csr_mtime_full[56]), .QN(n6876) );
  DFF_X1 pipeline_csr_mtime_full_reg_24_ ( .D(pipeline_csr_N2125), .CK(clk), 
        .Q(pipeline_csr_mtime_full[24]) );
  DFF_X1 pipeline_csr_time_full_reg_56_ ( .D(pipeline_csr_N2008), .CK(clk), 
        .Q(pipeline_csr_time_full[56]), .QN(n6877) );
  DFF_X1 pipeline_csr_time_full_reg_24_ ( .D(pipeline_csr_N1976), .CK(clk), 
        .Q(pipeline_csr_time_full[24]), .QN(n6833) );
  DFF_X1 pipeline_csr_cycle_full_reg_56_ ( .D(pipeline_csr_N1944), .CK(clk), 
        .Q(pipeline_csr_cycle_full[56]) );
  DFF_X1 pipeline_csr_cycle_full_reg_24_ ( .D(pipeline_csr_N1912), .CK(clk), 
        .Q(pipeline_csr_cycle_full[24]) );
  DFF_X1 pipeline_csr_mtime_full_reg_55_ ( .D(pipeline_csr_N2156), .CK(clk), 
        .Q(pipeline_csr_mtime_full[55]), .QN(n6878) );
  DFF_X1 pipeline_csr_mtime_full_reg_23_ ( .D(pipeline_csr_N2124), .CK(clk), 
        .Q(pipeline_csr_mtime_full[23]) );
  DFF_X1 pipeline_csr_time_full_reg_55_ ( .D(pipeline_csr_N2007), .CK(clk), 
        .Q(pipeline_csr_time_full[55]), .QN(n6879) );
  DFF_X1 pipeline_csr_time_full_reg_23_ ( .D(pipeline_csr_N1975), .CK(clk), 
        .Q(pipeline_csr_time_full[23]), .QN(n6900) );
  DFF_X1 pipeline_csr_cycle_full_reg_55_ ( .D(pipeline_csr_N1943), .CK(clk), 
        .Q(pipeline_csr_cycle_full[55]) );
  DFF_X1 pipeline_csr_cycle_full_reg_23_ ( .D(pipeline_csr_N1911), .CK(clk), 
        .Q(pipeline_csr_cycle_full[23]) );
  DFF_X1 pipeline_csr_mtime_full_reg_54_ ( .D(pipeline_csr_N2155), .CK(clk), 
        .Q(pipeline_csr_mtime_full[54]), .QN(n6910) );
  DFF_X1 pipeline_csr_mtime_full_reg_37_ ( .D(pipeline_csr_N2138), .CK(clk), 
        .Q(pipeline_csr_mtime_full[37]) );
  DFF_X1 pipeline_csr_mtime_full_reg_5_ ( .D(pipeline_csr_N2106), .CK(clk), 
        .Q(pipeline_csr_mtime_full[5]), .QN(n6751) );
  DFF_X1 pipeline_csr_time_full_reg_37_ ( .D(pipeline_csr_N1989), .CK(clk), 
        .Q(pipeline_csr_time_full[37]) );
  DFF_X1 pipeline_csr_time_full_reg_5_ ( .D(pipeline_csr_N1957), .CK(clk), .Q(
        pipeline_csr_time_full[5]), .QN(n6891) );
  DFF_X1 pipeline_csr_cycle_full_reg_37_ ( .D(pipeline_csr_N1925), .CK(clk), 
        .Q(pipeline_csr_cycle_full[37]) );
  DFF_X1 pipeline_csr_cycle_full_reg_5_ ( .D(pipeline_csr_N1893), .CK(clk), 
        .Q(pipeline_csr_cycle_full[5]), .QN(n6890) );
  DFF_X1 pipeline_csr_mbadaddr_reg_3_ ( .D(n5809), .CK(clk), .Q(
        pipeline_csr_mbadaddr[3]), .QN(n6923) );
  DFF_X1 pipeline_regfile_data_reg_1__3_ ( .D(n5466), .CK(clk), .Q(
        pipeline_regfile_data[35]) );
  DFF_X1 pipeline_regfile_data_reg_2__3_ ( .D(n5467), .CK(clk), .Q(
        pipeline_regfile_data[67]) );
  DFF_X1 pipeline_regfile_data_reg_3__3_ ( .D(n5468), .CK(clk), .Q(
        pipeline_regfile_data[99]) );
  DFF_X1 pipeline_regfile_data_reg_4__3_ ( .D(n5469), .CK(clk), .Q(
        pipeline_regfile_data[131]) );
  DFF_X1 pipeline_regfile_data_reg_5__3_ ( .D(n5470), .CK(clk), .Q(
        pipeline_regfile_data[163]) );
  DFF_X1 pipeline_regfile_data_reg_6__3_ ( .D(n5471), .CK(clk), .Q(
        pipeline_regfile_data[195]) );
  DFF_X1 pipeline_regfile_data_reg_7__3_ ( .D(n5472), .CK(clk), .Q(
        pipeline_regfile_data[227]) );
  DFF_X1 pipeline_regfile_data_reg_8__3_ ( .D(n5473), .CK(clk), .Q(
        pipeline_regfile_data[259]) );
  DFF_X1 pipeline_regfile_data_reg_9__3_ ( .D(n5474), .CK(clk), .Q(
        pipeline_regfile_data[291]) );
  DFF_X1 pipeline_regfile_data_reg_10__3_ ( .D(n5475), .CK(clk), .Q(
        pipeline_regfile_data[323]) );
  DFF_X1 pipeline_regfile_data_reg_11__3_ ( .D(n5476), .CK(clk), .Q(
        pipeline_regfile_data[355]) );
  DFF_X1 pipeline_regfile_data_reg_12__3_ ( .D(n5477), .CK(clk), .Q(
        pipeline_regfile_data[387]) );
  DFF_X1 pipeline_regfile_data_reg_13__3_ ( .D(n5478), .CK(clk), .Q(
        pipeline_regfile_data[419]) );
  DFF_X1 pipeline_regfile_data_reg_14__3_ ( .D(n5479), .CK(clk), .Q(
        pipeline_regfile_data[451]) );
  DFF_X1 pipeline_regfile_data_reg_15__3_ ( .D(n5480), .CK(clk), .Q(
        pipeline_regfile_data[483]) );
  DFF_X1 pipeline_regfile_data_reg_16__3_ ( .D(n5481), .CK(clk), .Q(
        pipeline_regfile_data[515]) );
  DFF_X1 pipeline_regfile_data_reg_18__3_ ( .D(n5483), .CK(clk), .Q(
        pipeline_regfile_data[579]) );
  DFF_X1 pipeline_regfile_data_reg_19__3_ ( .D(n5484), .CK(clk), .Q(
        pipeline_regfile_data[611]) );
  DFF_X1 pipeline_regfile_data_reg_20__3_ ( .D(n5485), .CK(clk), .Q(
        pipeline_regfile_data[643]) );
  DFF_X1 pipeline_regfile_data_reg_21__3_ ( .D(n5486), .CK(clk), .Q(
        pipeline_regfile_data[675]) );
  DFF_X1 pipeline_regfile_data_reg_22__3_ ( .D(n5487), .CK(clk), .Q(
        pipeline_regfile_data[707]) );
  DFF_X1 pipeline_regfile_data_reg_23__3_ ( .D(n5488), .CK(clk), .Q(
        pipeline_regfile_data[739]) );
  DFF_X1 pipeline_regfile_data_reg_24__3_ ( .D(n5489), .CK(clk), .Q(
        pipeline_regfile_data[771]) );
  DFF_X1 pipeline_regfile_data_reg_26__3_ ( .D(n5491), .CK(clk), .Q(
        pipeline_regfile_data[835]) );
  DFF_X1 pipeline_regfile_data_reg_27__3_ ( .D(n5492), .CK(clk), .Q(
        pipeline_regfile_data[867]) );
  DFF_X1 pipeline_regfile_data_reg_28__3_ ( .D(n5493), .CK(clk), .Q(
        pipeline_regfile_data[899]) );
  DFF_X1 pipeline_regfile_data_reg_29__3_ ( .D(n5494), .CK(clk), .Q(
        pipeline_regfile_data[931]) );
  DFF_X1 pipeline_regfile_data_reg_30__3_ ( .D(n5495), .CK(clk), .Q(
        pipeline_regfile_data[963]) );
  DFF_X1 pipeline_regfile_data_reg_31__3_ ( .D(n5496), .CK(clk), .Q(
        pipeline_regfile_data[995]) );
  DFF_X1 pipeline_regfile_data_reg_1__1_ ( .D(n5528), .CK(clk), .Q(
        pipeline_regfile_data[33]) );
  DFF_X1 pipeline_regfile_data_reg_2__1_ ( .D(n5529), .CK(clk), .Q(
        pipeline_regfile_data[65]) );
  DFF_X1 pipeline_regfile_data_reg_3__1_ ( .D(n5530), .CK(clk), .Q(
        pipeline_regfile_data[97]) );
  DFF_X1 pipeline_regfile_data_reg_4__1_ ( .D(n5531), .CK(clk), .Q(
        pipeline_regfile_data[129]) );
  DFF_X1 pipeline_regfile_data_reg_5__1_ ( .D(n5532), .CK(clk), .Q(
        pipeline_regfile_data[161]) );
  DFF_X1 pipeline_regfile_data_reg_6__1_ ( .D(n5533), .CK(clk), .Q(
        pipeline_regfile_data[193]) );
  DFF_X1 pipeline_regfile_data_reg_7__1_ ( .D(n5534), .CK(clk), .Q(
        pipeline_regfile_data[225]) );
  DFF_X1 pipeline_regfile_data_reg_8__1_ ( .D(n5535), .CK(clk), .Q(
        pipeline_regfile_data[257]) );
  DFF_X1 pipeline_regfile_data_reg_9__1_ ( .D(n5536), .CK(clk), .Q(
        pipeline_regfile_data[289]) );
  DFF_X1 pipeline_regfile_data_reg_10__1_ ( .D(n5537), .CK(clk), .Q(
        pipeline_regfile_data[321]) );
  DFF_X1 pipeline_regfile_data_reg_11__1_ ( .D(n5538), .CK(clk), .Q(
        pipeline_regfile_data[353]) );
  DFF_X1 pipeline_regfile_data_reg_12__1_ ( .D(n5539), .CK(clk), .Q(
        pipeline_regfile_data[385]) );
  DFF_X1 pipeline_regfile_data_reg_13__1_ ( .D(n5540), .CK(clk), .Q(
        pipeline_regfile_data[417]) );
  DFF_X1 pipeline_regfile_data_reg_14__1_ ( .D(n5541), .CK(clk), .Q(
        pipeline_regfile_data[449]) );
  DFF_X1 pipeline_regfile_data_reg_15__1_ ( .D(n5542), .CK(clk), .Q(
        pipeline_regfile_data[481]) );
  DFF_X1 pipeline_regfile_data_reg_16__1_ ( .D(n5543), .CK(clk), .Q(
        pipeline_regfile_data[513]) );
  DFF_X1 pipeline_regfile_data_reg_17__1_ ( .D(n5544), .CK(clk), .Q(
        pipeline_regfile_data[545]) );
  DFF_X1 pipeline_regfile_data_reg_18__1_ ( .D(n5545), .CK(clk), .Q(
        pipeline_regfile_data[577]) );
  DFF_X1 pipeline_regfile_data_reg_19__1_ ( .D(n5546), .CK(clk), .Q(
        pipeline_regfile_data[609]) );
  DFF_X1 pipeline_regfile_data_reg_20__1_ ( .D(n5547), .CK(clk), .Q(
        pipeline_regfile_data[641]) );
  DFF_X1 pipeline_regfile_data_reg_21__1_ ( .D(n5548), .CK(clk), .Q(
        pipeline_regfile_data[673]) );
  DFF_X1 pipeline_regfile_data_reg_22__1_ ( .D(n5549), .CK(clk), .Q(
        pipeline_regfile_data[705]) );
  DFF_X1 pipeline_regfile_data_reg_23__1_ ( .D(n5550), .CK(clk), .Q(
        pipeline_regfile_data[737]) );
  DFF_X1 pipeline_regfile_data_reg_24__1_ ( .D(n5551), .CK(clk), .Q(
        pipeline_regfile_data[769]) );
  DFF_X1 pipeline_regfile_data_reg_25__1_ ( .D(n5552), .CK(clk), .Q(
        pipeline_regfile_data[801]) );
  DFF_X1 pipeline_regfile_data_reg_26__1_ ( .D(n5553), .CK(clk), .Q(
        pipeline_regfile_data[833]) );
  DFF_X1 pipeline_regfile_data_reg_27__1_ ( .D(n5554), .CK(clk), .Q(
        pipeline_regfile_data[865]) );
  DFF_X1 pipeline_regfile_data_reg_28__1_ ( .D(n5555), .CK(clk), .Q(
        pipeline_regfile_data[897]) );
  DFF_X1 pipeline_regfile_data_reg_29__1_ ( .D(n5556), .CK(clk), .Q(
        pipeline_regfile_data[929]) );
  DFF_X1 pipeline_regfile_data_reg_30__1_ ( .D(n5557), .CK(clk), .Q(
        pipeline_regfile_data[961]) );
  DFF_X1 pipeline_regfile_data_reg_31__1_ ( .D(n5558), .CK(clk), .Q(
        pipeline_regfile_data[993]) );
  DFF_X1 pipeline_csr_mtime_full_reg_33_ ( .D(pipeline_csr_N2134), .CK(clk), 
        .Q(pipeline_csr_mtime_full[33]) );
  DFF_X1 pipeline_csr_mtime_full_reg_1_ ( .D(pipeline_csr_N2102), .CK(clk), 
        .Q(pipeline_csr_mtime_full[1]), .QN(n6815) );
  DFF_X1 pipeline_csr_time_full_reg_33_ ( .D(pipeline_csr_N1985), .CK(clk), 
        .Q(pipeline_csr_time_full[33]) );
  DFF_X1 pipeline_csr_time_full_reg_1_ ( .D(pipeline_csr_N1953), .CK(clk), .Q(
        pipeline_csr_time_full[1]) );
  DFF_X1 pipeline_csr_cycle_full_reg_33_ ( .D(pipeline_csr_N1921), .CK(clk), 
        .Q(pipeline_csr_cycle_full[33]), .QN(n6817) );
  DFF_X1 pipeline_csr_cycle_full_reg_1_ ( .D(pipeline_csr_N1889), .CK(clk), 
        .Q(pipeline_csr_cycle_full[1]) );
  DFF_X1 pipeline_regfile_data_reg_1__4_ ( .D(n5435), .CK(clk), .Q(
        pipeline_regfile_data[36]) );
  DFF_X1 pipeline_regfile_data_reg_2__4_ ( .D(n5436), .CK(clk), .Q(
        pipeline_regfile_data[68]) );
  DFF_X1 pipeline_regfile_data_reg_3__4_ ( .D(n5437), .CK(clk), .Q(
        pipeline_regfile_data[100]) );
  DFF_X1 pipeline_regfile_data_reg_4__4_ ( .D(n5438), .CK(clk), .Q(
        pipeline_regfile_data[132]) );
  DFF_X1 pipeline_regfile_data_reg_5__4_ ( .D(n5439), .CK(clk), .Q(
        pipeline_regfile_data[164]) );
  DFF_X1 pipeline_regfile_data_reg_6__4_ ( .D(n5440), .CK(clk), .Q(
        pipeline_regfile_data[196]) );
  DFF_X1 pipeline_regfile_data_reg_7__4_ ( .D(n5441), .CK(clk), .Q(
        pipeline_regfile_data[228]) );
  DFF_X1 pipeline_regfile_data_reg_8__4_ ( .D(n5442), .CK(clk), .Q(
        pipeline_regfile_data[260]) );
  DFF_X1 pipeline_regfile_data_reg_9__4_ ( .D(n5443), .CK(clk), .Q(
        pipeline_regfile_data[292]) );
  DFF_X1 pipeline_regfile_data_reg_10__4_ ( .D(n5444), .CK(clk), .Q(
        pipeline_regfile_data[324]) );
  DFF_X1 pipeline_regfile_data_reg_11__4_ ( .D(n5445), .CK(clk), .Q(
        pipeline_regfile_data[356]) );
  DFF_X1 pipeline_regfile_data_reg_12__4_ ( .D(n5446), .CK(clk), .Q(
        pipeline_regfile_data[388]) );
  DFF_X1 pipeline_regfile_data_reg_13__4_ ( .D(n5447), .CK(clk), .Q(
        pipeline_regfile_data[420]) );
  DFF_X1 pipeline_regfile_data_reg_14__4_ ( .D(n5448), .CK(clk), .Q(
        pipeline_regfile_data[452]) );
  DFF_X1 pipeline_regfile_data_reg_15__4_ ( .D(n5449), .CK(clk), .Q(
        pipeline_regfile_data[484]) );
  DFF_X1 pipeline_regfile_data_reg_16__4_ ( .D(n5450), .CK(clk), .Q(
        pipeline_regfile_data[516]) );
  DFF_X1 pipeline_regfile_data_reg_17__4_ ( .D(n5451), .CK(clk), .Q(
        pipeline_regfile_data[548]) );
  DFF_X1 pipeline_regfile_data_reg_18__4_ ( .D(n5452), .CK(clk), .Q(
        pipeline_regfile_data[580]) );
  DFF_X1 pipeline_regfile_data_reg_20__4_ ( .D(n5454), .CK(clk), .Q(
        pipeline_regfile_data[644]) );
  DFF_X1 pipeline_regfile_data_reg_21__4_ ( .D(n5455), .CK(clk), .Q(
        pipeline_regfile_data[676]) );
  DFF_X1 pipeline_regfile_data_reg_22__4_ ( .D(n5456), .CK(clk), .Q(
        pipeline_regfile_data[708]) );
  DFF_X1 pipeline_regfile_data_reg_23__4_ ( .D(n5457), .CK(clk), .Q(
        pipeline_regfile_data[740]) );
  DFF_X1 pipeline_regfile_data_reg_24__4_ ( .D(n5458), .CK(clk), .Q(
        pipeline_regfile_data[772]) );
  DFF_X1 pipeline_regfile_data_reg_25__4_ ( .D(n5459), .CK(clk), .Q(
        pipeline_regfile_data[804]) );
  DFF_X1 pipeline_regfile_data_reg_26__4_ ( .D(n5460), .CK(clk), .Q(
        pipeline_regfile_data[836]) );
  DFF_X1 pipeline_regfile_data_reg_27__4_ ( .D(n5461), .CK(clk), .Q(
        pipeline_regfile_data[868]) );
  DFF_X1 pipeline_regfile_data_reg_28__4_ ( .D(n5462), .CK(clk), .Q(
        pipeline_regfile_data[900]) );
  DFF_X1 pipeline_regfile_data_reg_29__4_ ( .D(n5463), .CK(clk), .Q(
        pipeline_regfile_data[932]) );
  DFF_X1 pipeline_regfile_data_reg_30__4_ ( .D(n5464), .CK(clk), .Q(
        pipeline_regfile_data[964]) );
  DFF_X1 pipeline_regfile_data_reg_31__4_ ( .D(n5465), .CK(clk), .Q(
        pipeline_regfile_data[996]) );
  DFF_X1 pipeline_csr_mtime_full_reg_36_ ( .D(pipeline_csr_N2137), .CK(clk), 
        .Q(pipeline_csr_mtime_full[36]) );
  DFF_X1 pipeline_csr_mtime_full_reg_4_ ( .D(pipeline_csr_N2105), .CK(clk), 
        .Q(pipeline_csr_mtime_full[4]), .QN(n6827) );
  DFF_X1 pipeline_csr_time_full_reg_36_ ( .D(pipeline_csr_N1988), .CK(clk), 
        .Q(pipeline_csr_time_full[36]), .QN(n6836) );
  DFF_X1 pipeline_csr_time_full_reg_4_ ( .D(pipeline_csr_N1956), .CK(clk), .Q(
        pipeline_csr_time_full[4]) );
  DFF_X1 pipeline_csr_cycle_full_reg_36_ ( .D(pipeline_csr_N1924), .CK(clk), 
        .Q(pipeline_csr_cycle_full[36]) );
  DFF_X1 pipeline_csr_cycle_full_reg_4_ ( .D(pipeline_csr_N1892), .CK(clk), 
        .Q(pipeline_csr_cycle_full[4]) );
  DFF_X1 pipeline_regfile_data_reg_1__2_ ( .D(n5497), .CK(clk), .Q(
        pipeline_regfile_data[34]) );
  DFF_X1 pipeline_regfile_data_reg_2__2_ ( .D(n5498), .CK(clk), .Q(
        pipeline_regfile_data[66]) );
  DFF_X1 pipeline_regfile_data_reg_3__2_ ( .D(n5499), .CK(clk), .Q(
        pipeline_regfile_data[98]) );
  DFF_X1 pipeline_regfile_data_reg_4__2_ ( .D(n5500), .CK(clk), .Q(
        pipeline_regfile_data[130]) );
  DFF_X1 pipeline_regfile_data_reg_5__2_ ( .D(n5501), .CK(clk), .Q(
        pipeline_regfile_data[162]) );
  DFF_X1 pipeline_regfile_data_reg_6__2_ ( .D(n5502), .CK(clk), .Q(
        pipeline_regfile_data[194]) );
  DFF_X1 pipeline_regfile_data_reg_7__2_ ( .D(n5503), .CK(clk), .Q(
        pipeline_regfile_data[226]) );
  DFF_X1 pipeline_regfile_data_reg_8__2_ ( .D(n5504), .CK(clk), .Q(
        pipeline_regfile_data[258]) );
  DFF_X1 pipeline_regfile_data_reg_9__2_ ( .D(n5505), .CK(clk), .Q(
        pipeline_regfile_data[290]) );
  DFF_X1 pipeline_regfile_data_reg_10__2_ ( .D(n5506), .CK(clk), .Q(
        pipeline_regfile_data[322]) );
  DFF_X1 pipeline_regfile_data_reg_11__2_ ( .D(n5507), .CK(clk), .Q(
        pipeline_regfile_data[354]) );
  DFF_X1 pipeline_regfile_data_reg_12__2_ ( .D(n5508), .CK(clk), .Q(
        pipeline_regfile_data[386]) );
  DFF_X1 pipeline_regfile_data_reg_13__2_ ( .D(n5509), .CK(clk), .Q(
        pipeline_regfile_data[418]) );
  DFF_X1 pipeline_regfile_data_reg_14__2_ ( .D(n5510), .CK(clk), .Q(
        pipeline_regfile_data[450]) );
  DFF_X1 pipeline_regfile_data_reg_15__2_ ( .D(n5511), .CK(clk), .Q(
        pipeline_regfile_data[482]) );
  DFF_X1 pipeline_regfile_data_reg_16__2_ ( .D(n5512), .CK(clk), .Q(
        pipeline_regfile_data[514]) );
  DFF_X1 pipeline_regfile_data_reg_17__2_ ( .D(n5513), .CK(clk), .Q(
        pipeline_regfile_data[546]) );
  DFF_X1 pipeline_regfile_data_reg_18__2_ ( .D(n5514), .CK(clk), .Q(
        pipeline_regfile_data[578]) );
  DFF_X1 pipeline_regfile_data_reg_19__2_ ( .D(n5515), .CK(clk), .Q(
        pipeline_regfile_data[610]) );
  DFF_X1 pipeline_regfile_data_reg_20__2_ ( .D(n5516), .CK(clk), .Q(
        pipeline_regfile_data[642]) );
  DFF_X1 pipeline_regfile_data_reg_21__2_ ( .D(n5517), .CK(clk), .Q(
        pipeline_regfile_data[674]) );
  DFF_X1 pipeline_regfile_data_reg_22__2_ ( .D(n5518), .CK(clk), .Q(
        pipeline_regfile_data[706]) );
  DFF_X1 pipeline_regfile_data_reg_23__2_ ( .D(n5519), .CK(clk), .Q(
        pipeline_regfile_data[738]) );
  DFF_X1 pipeline_regfile_data_reg_24__2_ ( .D(n5520), .CK(clk), .Q(
        pipeline_regfile_data[770]) );
  DFF_X1 pipeline_regfile_data_reg_25__2_ ( .D(n5521), .CK(clk), .Q(
        pipeline_regfile_data[802]) );
  DFF_X1 pipeline_regfile_data_reg_26__2_ ( .D(n5522), .CK(clk), .Q(
        pipeline_regfile_data[834]) );
  DFF_X1 pipeline_regfile_data_reg_27__2_ ( .D(n5523), .CK(clk), .Q(
        pipeline_regfile_data[866]) );
  DFF_X1 pipeline_regfile_data_reg_28__2_ ( .D(n5524), .CK(clk), .Q(
        pipeline_regfile_data[898]) );
  DFF_X1 pipeline_regfile_data_reg_29__2_ ( .D(n5525), .CK(clk), .Q(
        pipeline_regfile_data[930]) );
  DFF_X1 pipeline_regfile_data_reg_30__2_ ( .D(n5526), .CK(clk), .Q(
        pipeline_regfile_data[962]) );
  DFF_X1 pipeline_regfile_data_reg_31__2_ ( .D(n5527), .CK(clk), .Q(
        pipeline_regfile_data[994]) );
  DFF_X1 pipeline_csr_mtime_full_reg_34_ ( .D(pipeline_csr_N2135), .CK(clk), 
        .Q(pipeline_csr_mtime_full[34]) );
  DFF_X1 pipeline_csr_mtime_full_reg_2_ ( .D(pipeline_csr_N2103), .CK(clk), 
        .Q(pipeline_csr_mtime_full[2]), .QN(n6850) );
  DFF_X1 pipeline_csr_time_full_reg_34_ ( .D(pipeline_csr_N1986), .CK(clk), 
        .Q(pipeline_csr_time_full[34]), .QN(n6835) );
  DFF_X1 pipeline_csr_time_full_reg_2_ ( .D(pipeline_csr_N1954), .CK(clk), .Q(
        pipeline_csr_time_full[2]) );
  DFF_X1 pipeline_csr_cycle_full_reg_34_ ( .D(pipeline_csr_N1922), .CK(clk), 
        .Q(pipeline_csr_cycle_full[34]) );
  DFF_X1 pipeline_csr_cycle_full_reg_2_ ( .D(pipeline_csr_N1890), .CK(clk), 
        .Q(pipeline_csr_cycle_full[2]) );
  DFF_X1 pipeline_regfile_data_reg_1__5_ ( .D(n5404), .CK(clk), .Q(
        pipeline_regfile_data[37]) );
  DFF_X1 pipeline_regfile_data_reg_2__5_ ( .D(n5405), .CK(clk), .Q(
        pipeline_regfile_data[69]) );
  DFF_X1 pipeline_regfile_data_reg_3__5_ ( .D(n5406), .CK(clk), .Q(
        pipeline_regfile_data[101]) );
  DFF_X1 pipeline_regfile_data_reg_4__5_ ( .D(n5407), .CK(clk), .Q(
        pipeline_regfile_data[133]) );
  DFF_X1 pipeline_regfile_data_reg_5__5_ ( .D(n5408), .CK(clk), .Q(
        pipeline_regfile_data[165]) );
  DFF_X1 pipeline_regfile_data_reg_6__5_ ( .D(n5409), .CK(clk), .Q(
        pipeline_regfile_data[197]) );
  DFF_X1 pipeline_regfile_data_reg_7__5_ ( .D(n5410), .CK(clk), .Q(
        pipeline_regfile_data[229]) );
  DFF_X1 pipeline_regfile_data_reg_8__5_ ( .D(n5411), .CK(clk), .Q(
        pipeline_regfile_data[261]) );
  DFF_X1 pipeline_regfile_data_reg_9__5_ ( .D(n5412), .CK(clk), .Q(
        pipeline_regfile_data[293]) );
  DFF_X1 pipeline_regfile_data_reg_10__5_ ( .D(n5413), .CK(clk), .Q(
        pipeline_regfile_data[325]) );
  DFF_X1 pipeline_regfile_data_reg_11__5_ ( .D(n5414), .CK(clk), .Q(
        pipeline_regfile_data[357]) );
  DFF_X1 pipeline_regfile_data_reg_12__5_ ( .D(n5415), .CK(clk), .Q(
        pipeline_regfile_data[389]) );
  DFF_X1 pipeline_regfile_data_reg_13__5_ ( .D(n5416), .CK(clk), .Q(
        pipeline_regfile_data[421]) );
  DFF_X1 pipeline_regfile_data_reg_14__5_ ( .D(n5417), .CK(clk), .Q(
        pipeline_regfile_data[453]) );
  DFF_X1 pipeline_regfile_data_reg_15__5_ ( .D(n5418), .CK(clk), .Q(
        pipeline_regfile_data[485]) );
  DFF_X1 pipeline_regfile_data_reg_16__5_ ( .D(n5419), .CK(clk), .Q(
        pipeline_regfile_data[517]) );
  DFF_X1 pipeline_regfile_data_reg_17__5_ ( .D(n5420), .CK(clk), .Q(
        pipeline_regfile_data[549]) );
  DFF_X1 pipeline_regfile_data_reg_18__5_ ( .D(n5421), .CK(clk), .Q(
        pipeline_regfile_data[581]) );
  DFF_X1 pipeline_regfile_data_reg_19__5_ ( .D(n5422), .CK(clk), .Q(
        pipeline_regfile_data[613]) );
  DFF_X1 pipeline_regfile_data_reg_20__5_ ( .D(n5423), .CK(clk), .Q(
        pipeline_regfile_data[645]) );
  DFF_X1 pipeline_regfile_data_reg_21__5_ ( .D(n5424), .CK(clk), .Q(
        pipeline_regfile_data[677]) );
  DFF_X1 pipeline_regfile_data_reg_22__5_ ( .D(n5425), .CK(clk), .Q(
        pipeline_regfile_data[709]) );
  DFF_X1 pipeline_regfile_data_reg_23__5_ ( .D(n5426), .CK(clk), .Q(
        pipeline_regfile_data[741]) );
  DFF_X1 pipeline_regfile_data_reg_24__5_ ( .D(n5427), .CK(clk), .Q(
        pipeline_regfile_data[773]) );
  DFF_X1 pipeline_regfile_data_reg_25__5_ ( .D(n5428), .CK(clk), .Q(
        pipeline_regfile_data[805]) );
  DFF_X1 pipeline_regfile_data_reg_26__5_ ( .D(n5429), .CK(clk), .Q(
        pipeline_regfile_data[837]) );
  DFF_X1 pipeline_regfile_data_reg_27__5_ ( .D(n5430), .CK(clk), .Q(
        pipeline_regfile_data[869]) );
  DFF_X1 pipeline_regfile_data_reg_28__5_ ( .D(n5431), .CK(clk), .Q(
        pipeline_regfile_data[901]) );
  DFF_X1 pipeline_regfile_data_reg_29__5_ ( .D(n5432), .CK(clk), .Q(
        pipeline_regfile_data[933]) );
  DFF_X1 pipeline_regfile_data_reg_30__5_ ( .D(n5433), .CK(clk), .Q(
        pipeline_regfile_data[965]) );
  DFF_X1 pipeline_regfile_data_reg_31__5_ ( .D(n5434), .CK(clk), .Q(
        pipeline_regfile_data[997]) );
  DFF_X1 pipeline_csr_mtime_full_reg_38_ ( .D(pipeline_csr_N2139), .CK(clk), 
        .Q(pipeline_csr_mtime_full[38]) );
  DFF_X2 pipeline_csr_instret_full_reg_6_ ( .D(n6040), .CK(clk), .Q(
        pipeline_csr_instret_full[6]), .QN(n1389) );
  DFF_X1 pipeline_csr_mtime_full_reg_6_ ( .D(pipeline_csr_N2107), .CK(clk), 
        .Q(pipeline_csr_mtime_full[6]), .QN(n6824) );
  DFF_X1 pipeline_csr_time_full_reg_38_ ( .D(pipeline_csr_N1990), .CK(clk), 
        .Q(pipeline_csr_time_full[38]), .QN(n6913) );
  DFF_X1 pipeline_csr_time_full_reg_6_ ( .D(pipeline_csr_N1958), .CK(clk), .Q(
        pipeline_csr_time_full[6]) );
  DFF_X2 pipeline_csr_cycle_full_reg_38_ ( .D(pipeline_csr_N1926), .CK(clk), 
        .Q(pipeline_csr_cycle_full[38]), .QN(n1160) );
  DFF_X1 pipeline_csr_cycle_full_reg_6_ ( .D(pipeline_csr_N1894), .CK(clk), 
        .Q(pipeline_csr_cycle_full[6]) );
  DFF_X1 pipeline_regfile_data_reg_1__6_ ( .D(n5373), .CK(clk), .Q(
        pipeline_regfile_data[38]) );
  DFF_X1 pipeline_regfile_data_reg_2__6_ ( .D(n5374), .CK(clk), .Q(
        pipeline_regfile_data[70]) );
  DFF_X1 pipeline_regfile_data_reg_3__6_ ( .D(n5375), .CK(clk), .Q(
        pipeline_regfile_data[102]) );
  DFF_X1 pipeline_regfile_data_reg_4__6_ ( .D(n5376), .CK(clk), .Q(
        pipeline_regfile_data[134]) );
  DFF_X1 pipeline_regfile_data_reg_5__6_ ( .D(n5377), .CK(clk), .Q(
        pipeline_regfile_data[166]) );
  DFF_X1 pipeline_regfile_data_reg_6__6_ ( .D(n5378), .CK(clk), .Q(
        pipeline_regfile_data[198]) );
  DFF_X1 pipeline_regfile_data_reg_7__6_ ( .D(n5379), .CK(clk), .Q(
        pipeline_regfile_data[230]) );
  DFF_X1 pipeline_regfile_data_reg_8__6_ ( .D(n5380), .CK(clk), .Q(
        pipeline_regfile_data[262]) );
  DFF_X1 pipeline_regfile_data_reg_9__6_ ( .D(n5381), .CK(clk), .Q(
        pipeline_regfile_data[294]) );
  DFF_X1 pipeline_regfile_data_reg_10__6_ ( .D(n5382), .CK(clk), .Q(
        pipeline_regfile_data[326]) );
  DFF_X1 pipeline_regfile_data_reg_11__6_ ( .D(n5383), .CK(clk), .Q(
        pipeline_regfile_data[358]) );
  DFF_X1 pipeline_regfile_data_reg_12__6_ ( .D(n5384), .CK(clk), .Q(
        pipeline_regfile_data[390]) );
  DFF_X1 pipeline_regfile_data_reg_13__6_ ( .D(n5385), .CK(clk), .Q(
        pipeline_regfile_data[422]) );
  DFF_X1 pipeline_regfile_data_reg_14__6_ ( .D(n5386), .CK(clk), .Q(
        pipeline_regfile_data[454]) );
  DFF_X1 pipeline_regfile_data_reg_15__6_ ( .D(n5387), .CK(clk), .Q(
        pipeline_regfile_data[486]) );
  DFF_X1 pipeline_regfile_data_reg_16__6_ ( .D(n5388), .CK(clk), .Q(
        pipeline_regfile_data[518]) );
  DFF_X1 pipeline_regfile_data_reg_17__6_ ( .D(n5389), .CK(clk), .Q(
        pipeline_regfile_data[550]) );
  DFF_X1 pipeline_regfile_data_reg_18__6_ ( .D(n5390), .CK(clk), .Q(
        pipeline_regfile_data[582]) );
  DFF_X1 pipeline_regfile_data_reg_19__6_ ( .D(n5391), .CK(clk), .Q(
        pipeline_regfile_data[614]) );
  DFF_X1 pipeline_regfile_data_reg_20__6_ ( .D(n5392), .CK(clk), .Q(
        pipeline_regfile_data[646]) );
  DFF_X1 pipeline_regfile_data_reg_21__6_ ( .D(n5393), .CK(clk), .Q(
        pipeline_regfile_data[678]) );
  DFF_X1 pipeline_regfile_data_reg_22__6_ ( .D(n5394), .CK(clk), .Q(
        pipeline_regfile_data[710]) );
  DFF_X1 pipeline_regfile_data_reg_23__6_ ( .D(n5395), .CK(clk), .Q(
        pipeline_regfile_data[742]) );
  DFF_X1 pipeline_regfile_data_reg_24__6_ ( .D(n5396), .CK(clk), .Q(
        pipeline_regfile_data[774]) );
  DFF_X1 pipeline_regfile_data_reg_25__6_ ( .D(n5397), .CK(clk), .Q(
        pipeline_regfile_data[806]) );
  DFF_X1 pipeline_regfile_data_reg_26__6_ ( .D(n5398), .CK(clk), .Q(
        pipeline_regfile_data[838]) );
  DFF_X1 pipeline_regfile_data_reg_27__6_ ( .D(n5399), .CK(clk), .Q(
        pipeline_regfile_data[870]) );
  DFF_X1 pipeline_regfile_data_reg_28__6_ ( .D(n5400), .CK(clk), .Q(
        pipeline_regfile_data[902]) );
  DFF_X1 pipeline_regfile_data_reg_29__6_ ( .D(n5401), .CK(clk), .Q(
        pipeline_regfile_data[934]) );
  DFF_X1 pipeline_regfile_data_reg_30__6_ ( .D(n5402), .CK(clk), .Q(
        pipeline_regfile_data[966]) );
  DFF_X1 pipeline_regfile_data_reg_31__6_ ( .D(n5403), .CK(clk), .Q(
        pipeline_regfile_data[998]) );
  DFF_X1 pipeline_regfile_data_reg_1__7_ ( .D(n5342), .CK(clk), .Q(
        pipeline_regfile_data[39]) );
  DFF_X1 pipeline_regfile_data_reg_2__7_ ( .D(n5343), .CK(clk), .Q(
        pipeline_regfile_data[71]) );
  DFF_X1 pipeline_regfile_data_reg_3__7_ ( .D(n5344), .CK(clk), .Q(
        pipeline_regfile_data[103]) );
  DFF_X1 pipeline_regfile_data_reg_4__7_ ( .D(n5345), .CK(clk), .Q(
        pipeline_regfile_data[135]) );
  DFF_X1 pipeline_regfile_data_reg_5__7_ ( .D(n5346), .CK(clk), .Q(
        pipeline_regfile_data[167]) );
  DFF_X1 pipeline_regfile_data_reg_6__7_ ( .D(n5347), .CK(clk), .Q(
        pipeline_regfile_data[199]) );
  DFF_X1 pipeline_regfile_data_reg_7__7_ ( .D(n5348), .CK(clk), .Q(
        pipeline_regfile_data[231]) );
  DFF_X1 pipeline_regfile_data_reg_8__7_ ( .D(n5349), .CK(clk), .Q(
        pipeline_regfile_data[263]) );
  DFF_X1 pipeline_regfile_data_reg_9__7_ ( .D(n5350), .CK(clk), .Q(
        pipeline_regfile_data[295]) );
  DFF_X1 pipeline_regfile_data_reg_10__7_ ( .D(n5351), .CK(clk), .Q(
        pipeline_regfile_data[327]) );
  DFF_X1 pipeline_regfile_data_reg_11__7_ ( .D(n5352), .CK(clk), .Q(
        pipeline_regfile_data[359]) );
  DFF_X1 pipeline_regfile_data_reg_12__7_ ( .D(n5353), .CK(clk), .Q(
        pipeline_regfile_data[391]) );
  DFF_X1 pipeline_regfile_data_reg_13__7_ ( .D(n5354), .CK(clk), .Q(
        pipeline_regfile_data[423]) );
  DFF_X1 pipeline_regfile_data_reg_14__7_ ( .D(n5355), .CK(clk), .Q(
        pipeline_regfile_data[455]) );
  DFF_X1 pipeline_regfile_data_reg_15__7_ ( .D(n5356), .CK(clk), .Q(
        pipeline_regfile_data[487]) );
  DFF_X1 pipeline_regfile_data_reg_16__7_ ( .D(n5357), .CK(clk), .Q(
        pipeline_regfile_data[519]) );
  DFF_X1 pipeline_regfile_data_reg_17__7_ ( .D(n5358), .CK(clk), .Q(
        pipeline_regfile_data[551]) );
  DFF_X1 pipeline_regfile_data_reg_18__7_ ( .D(n5359), .CK(clk), .Q(
        pipeline_regfile_data[583]) );
  DFF_X1 pipeline_regfile_data_reg_19__7_ ( .D(n5360), .CK(clk), .Q(
        pipeline_regfile_data[615]) );
  DFF_X1 pipeline_regfile_data_reg_20__7_ ( .D(n5361), .CK(clk), .Q(
        pipeline_regfile_data[647]) );
  DFF_X1 pipeline_regfile_data_reg_21__7_ ( .D(n5362), .CK(clk), .Q(
        pipeline_regfile_data[679]) );
  DFF_X1 pipeline_regfile_data_reg_22__7_ ( .D(n5363), .CK(clk), .Q(
        pipeline_regfile_data[711]) );
  DFF_X1 pipeline_regfile_data_reg_23__7_ ( .D(n5364), .CK(clk), .Q(
        pipeline_regfile_data[743]) );
  DFF_X1 pipeline_regfile_data_reg_24__7_ ( .D(n5365), .CK(clk), .Q(
        pipeline_regfile_data[775]) );
  DFF_X1 pipeline_regfile_data_reg_25__7_ ( .D(n5366), .CK(clk), .Q(
        pipeline_regfile_data[807]) );
  DFF_X1 pipeline_regfile_data_reg_26__7_ ( .D(n5367), .CK(clk), .Q(
        pipeline_regfile_data[839]) );
  DFF_X1 pipeline_regfile_data_reg_27__7_ ( .D(n5368), .CK(clk), .Q(
        pipeline_regfile_data[871]) );
  DFF_X1 pipeline_regfile_data_reg_28__7_ ( .D(n5369), .CK(clk), .Q(
        pipeline_regfile_data[903]) );
  DFF_X1 pipeline_regfile_data_reg_29__7_ ( .D(n5370), .CK(clk), .Q(
        pipeline_regfile_data[935]) );
  DFF_X1 pipeline_regfile_data_reg_30__7_ ( .D(n5371), .CK(clk), .Q(
        pipeline_regfile_data[967]) );
  DFF_X1 pipeline_regfile_data_reg_31__7_ ( .D(n5372), .CK(clk), .Q(
        pipeline_regfile_data[999]) );
  DFF_X1 pipeline_csr_mtime_full_reg_40_ ( .D(pipeline_csr_N2141), .CK(clk), 
        .Q(pipeline_csr_mtime_full[40]) );
  DFF_X2 pipeline_csr_instret_full_reg_40_ ( .D(n6006), .CK(clk), .Q(n10618), 
        .QN(n1423) );
  DFF_X2 pipeline_csr_mtvec_reg_8_ ( .D(n6200), .CK(clk), .Q(n10635) );
  DFF_X1 pipeline_csr_mtime_full_reg_8_ ( .D(pipeline_csr_N2109), .CK(clk), 
        .Q(pipeline_csr_mtime_full[8]), .QN(n6825) );
  DFF_X2 pipeline_csr_time_full_reg_40_ ( .D(pipeline_csr_N1992), .CK(clk), 
        .Q(pipeline_csr_time_full[40]), .QN(n1157) );
  DFF_X1 pipeline_csr_time_full_reg_8_ ( .D(pipeline_csr_N1960), .CK(clk), .Q(
        pipeline_csr_time_full[8]) );
  DFF_X1 pipeline_csr_cycle_full_reg_40_ ( .D(pipeline_csr_N1928), .CK(clk), 
        .Q(pipeline_csr_cycle_full[40]), .QN(n6840) );
  DFF_X1 pipeline_csr_cycle_full_reg_8_ ( .D(pipeline_csr_N1896), .CK(clk), 
        .Q(pipeline_csr_cycle_full[8]) );
  DFF_X1 pipeline_regfile_data_reg_1__8_ ( .D(n5311), .CK(clk), .Q(
        pipeline_regfile_data[40]) );
  DFF_X1 pipeline_regfile_data_reg_2__8_ ( .D(n5312), .CK(clk), .Q(
        pipeline_regfile_data[72]) );
  DFF_X1 pipeline_regfile_data_reg_3__8_ ( .D(n5313), .CK(clk), .Q(
        pipeline_regfile_data[104]) );
  DFF_X1 pipeline_regfile_data_reg_4__8_ ( .D(n5314), .CK(clk), .Q(
        pipeline_regfile_data[136]) );
  DFF_X1 pipeline_regfile_data_reg_5__8_ ( .D(n5315), .CK(clk), .Q(
        pipeline_regfile_data[168]) );
  DFF_X1 pipeline_regfile_data_reg_6__8_ ( .D(n5316), .CK(clk), .Q(
        pipeline_regfile_data[200]) );
  DFF_X1 pipeline_regfile_data_reg_7__8_ ( .D(n5317), .CK(clk), .Q(
        pipeline_regfile_data[232]) );
  DFF_X1 pipeline_regfile_data_reg_8__8_ ( .D(n5318), .CK(clk), .Q(
        pipeline_regfile_data[264]) );
  DFF_X1 pipeline_regfile_data_reg_9__8_ ( .D(n5319), .CK(clk), .Q(
        pipeline_regfile_data[296]) );
  DFF_X1 pipeline_regfile_data_reg_10__8_ ( .D(n5320), .CK(clk), .Q(
        pipeline_regfile_data[328]) );
  DFF_X1 pipeline_regfile_data_reg_11__8_ ( .D(n5321), .CK(clk), .Q(
        pipeline_regfile_data[360]) );
  DFF_X1 pipeline_regfile_data_reg_12__8_ ( .D(n5322), .CK(clk), .Q(
        pipeline_regfile_data[392]) );
  DFF_X1 pipeline_regfile_data_reg_13__8_ ( .D(n5323), .CK(clk), .Q(
        pipeline_regfile_data[424]) );
  DFF_X1 pipeline_regfile_data_reg_14__8_ ( .D(n5324), .CK(clk), .Q(
        pipeline_regfile_data[456]) );
  DFF_X1 pipeline_regfile_data_reg_15__8_ ( .D(n5325), .CK(clk), .Q(
        pipeline_regfile_data[488]) );
  DFF_X1 pipeline_regfile_data_reg_16__8_ ( .D(n5326), .CK(clk), .Q(
        pipeline_regfile_data[520]) );
  DFF_X1 pipeline_regfile_data_reg_17__8_ ( .D(n5327), .CK(clk), .Q(
        pipeline_regfile_data[552]) );
  DFF_X1 pipeline_regfile_data_reg_18__8_ ( .D(n5328), .CK(clk), .Q(
        pipeline_regfile_data[584]) );
  DFF_X1 pipeline_regfile_data_reg_19__8_ ( .D(n5329), .CK(clk), .Q(
        pipeline_regfile_data[616]) );
  DFF_X1 pipeline_regfile_data_reg_20__8_ ( .D(n5330), .CK(clk), .Q(
        pipeline_regfile_data[648]) );
  DFF_X1 pipeline_regfile_data_reg_21__8_ ( .D(n5331), .CK(clk), .Q(
        pipeline_regfile_data[680]) );
  DFF_X1 pipeline_regfile_data_reg_22__8_ ( .D(n5332), .CK(clk), .Q(
        pipeline_regfile_data[712]) );
  DFF_X1 pipeline_regfile_data_reg_23__8_ ( .D(n5333), .CK(clk), .Q(
        pipeline_regfile_data[744]) );
  DFF_X1 pipeline_regfile_data_reg_24__8_ ( .D(n5334), .CK(clk), .Q(
        pipeline_regfile_data[776]) );
  DFF_X1 pipeline_regfile_data_reg_25__8_ ( .D(n5335), .CK(clk), .Q(
        pipeline_regfile_data[808]) );
  DFF_X1 pipeline_regfile_data_reg_26__8_ ( .D(n5336), .CK(clk), .Q(
        pipeline_regfile_data[840]) );
  DFF_X1 pipeline_regfile_data_reg_27__8_ ( .D(n5337), .CK(clk), .Q(
        pipeline_regfile_data[872]) );
  DFF_X1 pipeline_regfile_data_reg_28__8_ ( .D(n5338), .CK(clk), .Q(
        pipeline_regfile_data[904]) );
  DFF_X1 pipeline_regfile_data_reg_29__8_ ( .D(n5339), .CK(clk), .Q(
        pipeline_regfile_data[936]) );
  DFF_X1 pipeline_regfile_data_reg_30__8_ ( .D(n5340), .CK(clk), .Q(
        pipeline_regfile_data[968]) );
  DFF_X1 pipeline_regfile_data_reg_31__8_ ( .D(n5341), .CK(clk), .Q(
        pipeline_regfile_data[1000]) );
  DFF_X1 pipeline_csr_mtime_full_reg_41_ ( .D(pipeline_csr_N2142), .CK(clk), 
        .Q(pipeline_csr_mtime_full[41]), .QN(n6888) );
  DFF_X1 pipeline_csr_mtime_full_reg_9_ ( .D(pipeline_csr_N2110), .CK(clk), 
        .Q(pipeline_csr_mtime_full[9]), .QN(n6860) );
  DFF_X1 pipeline_csr_time_full_reg_41_ ( .D(pipeline_csr_N1993), .CK(clk), 
        .Q(pipeline_csr_time_full[41]) );
  DFF_X1 pipeline_csr_time_full_reg_9_ ( .D(pipeline_csr_N1961), .CK(clk), .Q(
        pipeline_csr_time_full[9]), .QN(n6889) );
  DFF_X1 pipeline_csr_cycle_full_reg_41_ ( .D(pipeline_csr_N1929), .CK(clk), 
        .Q(pipeline_csr_cycle_full[41]) );
  DFF_X1 pipeline_csr_cycle_full_reg_9_ ( .D(pipeline_csr_N1897), .CK(clk), 
        .Q(pipeline_csr_cycle_full[9]) );
  DFF_X1 pipeline_regfile_data_reg_1__9_ ( .D(n5280), .CK(clk), .Q(
        pipeline_regfile_data[41]) );
  DFF_X1 pipeline_regfile_data_reg_2__9_ ( .D(n5281), .CK(clk), .Q(
        pipeline_regfile_data[73]) );
  DFF_X1 pipeline_regfile_data_reg_3__9_ ( .D(n5282), .CK(clk), .Q(
        pipeline_regfile_data[105]) );
  DFF_X1 pipeline_regfile_data_reg_4__9_ ( .D(n5283), .CK(clk), .Q(
        pipeline_regfile_data[137]) );
  DFF_X1 pipeline_regfile_data_reg_5__9_ ( .D(n5284), .CK(clk), .Q(
        pipeline_regfile_data[169]) );
  DFF_X1 pipeline_regfile_data_reg_6__9_ ( .D(n5285), .CK(clk), .Q(
        pipeline_regfile_data[201]) );
  DFF_X1 pipeline_regfile_data_reg_7__9_ ( .D(n5286), .CK(clk), .Q(
        pipeline_regfile_data[233]) );
  DFF_X1 pipeline_regfile_data_reg_8__9_ ( .D(n5287), .CK(clk), .Q(
        pipeline_regfile_data[265]) );
  DFF_X1 pipeline_regfile_data_reg_9__9_ ( .D(n5288), .CK(clk), .Q(
        pipeline_regfile_data[297]) );
  DFF_X1 pipeline_regfile_data_reg_10__9_ ( .D(n5289), .CK(clk), .Q(
        pipeline_regfile_data[329]) );
  DFF_X1 pipeline_regfile_data_reg_11__9_ ( .D(n5290), .CK(clk), .Q(
        pipeline_regfile_data[361]) );
  DFF_X1 pipeline_regfile_data_reg_12__9_ ( .D(n5291), .CK(clk), .Q(
        pipeline_regfile_data[393]) );
  DFF_X1 pipeline_regfile_data_reg_13__9_ ( .D(n5292), .CK(clk), .Q(
        pipeline_regfile_data[425]) );
  DFF_X1 pipeline_regfile_data_reg_14__9_ ( .D(n5293), .CK(clk), .Q(
        pipeline_regfile_data[457]) );
  DFF_X1 pipeline_regfile_data_reg_15__9_ ( .D(n5294), .CK(clk), .Q(
        pipeline_regfile_data[489]) );
  DFF_X1 pipeline_regfile_data_reg_16__9_ ( .D(n5295), .CK(clk), .Q(
        pipeline_regfile_data[521]) );
  DFF_X1 pipeline_regfile_data_reg_17__9_ ( .D(n5296), .CK(clk), .Q(
        pipeline_regfile_data[553]) );
  DFF_X1 pipeline_regfile_data_reg_18__9_ ( .D(n5297), .CK(clk), .Q(
        pipeline_regfile_data[585]) );
  DFF_X1 pipeline_regfile_data_reg_19__9_ ( .D(n5298), .CK(clk), .Q(
        pipeline_regfile_data[617]) );
  DFF_X1 pipeline_regfile_data_reg_20__9_ ( .D(n5299), .CK(clk), .Q(
        pipeline_regfile_data[649]) );
  DFF_X1 pipeline_regfile_data_reg_21__9_ ( .D(n5300), .CK(clk), .Q(
        pipeline_regfile_data[681]) );
  DFF_X1 pipeline_regfile_data_reg_22__9_ ( .D(n5301), .CK(clk), .Q(
        pipeline_regfile_data[713]) );
  DFF_X1 pipeline_regfile_data_reg_23__9_ ( .D(n5302), .CK(clk), .Q(
        pipeline_regfile_data[745]) );
  DFF_X1 pipeline_regfile_data_reg_24__9_ ( .D(n5303), .CK(clk), .Q(
        pipeline_regfile_data[777]) );
  DFF_X1 pipeline_regfile_data_reg_25__9_ ( .D(n5304), .CK(clk), .Q(
        pipeline_regfile_data[809]) );
  DFF_X1 pipeline_regfile_data_reg_26__9_ ( .D(n5305), .CK(clk), .Q(
        pipeline_regfile_data[841]) );
  DFF_X1 pipeline_regfile_data_reg_27__9_ ( .D(n5306), .CK(clk), .Q(
        pipeline_regfile_data[873]) );
  DFF_X1 pipeline_regfile_data_reg_28__9_ ( .D(n5307), .CK(clk), .Q(
        pipeline_regfile_data[905]) );
  DFF_X1 pipeline_regfile_data_reg_29__9_ ( .D(n5308), .CK(clk), .Q(
        pipeline_regfile_data[937]) );
  DFF_X1 pipeline_regfile_data_reg_30__9_ ( .D(n5309), .CK(clk), .Q(
        pipeline_regfile_data[969]) );
  DFF_X1 pipeline_regfile_data_reg_31__9_ ( .D(n5310), .CK(clk), .Q(
        pipeline_regfile_data[1001]) );
  DFF_X1 pipeline_csr_mtime_full_reg_42_ ( .D(pipeline_csr_N2143), .CK(clk), 
        .Q(pipeline_csr_mtime_full[42]), .QN(n6908) );
  DFF_X1 pipeline_csr_mtime_full_reg_10_ ( .D(pipeline_csr_N2111), .CK(clk), 
        .Q(pipeline_csr_mtime_full[10]) );
  DFF_X1 pipeline_csr_time_full_reg_42_ ( .D(pipeline_csr_N1994), .CK(clk), 
        .Q(pipeline_csr_time_full[42]) );
  DFF_X1 pipeline_csr_time_full_reg_10_ ( .D(pipeline_csr_N1962), .CK(clk), 
        .Q(pipeline_csr_time_full[10]), .QN(n6884) );
  DFF_X1 pipeline_csr_cycle_full_reg_42_ ( .D(pipeline_csr_N1930), .CK(clk), 
        .Q(pipeline_csr_cycle_full[42]) );
  DFF_X1 pipeline_csr_cycle_full_reg_10_ ( .D(pipeline_csr_N1898), .CK(clk), 
        .Q(pipeline_csr_cycle_full[10]) );
  DFF_X1 pipeline_regfile_data_reg_1__10_ ( .D(n5249), .CK(clk), .Q(
        pipeline_regfile_data[42]) );
  DFF_X1 pipeline_regfile_data_reg_2__10_ ( .D(n5250), .CK(clk), .Q(
        pipeline_regfile_data[74]) );
  DFF_X1 pipeline_regfile_data_reg_3__10_ ( .D(n5251), .CK(clk), .Q(
        pipeline_regfile_data[106]) );
  DFF_X1 pipeline_regfile_data_reg_4__10_ ( .D(n5252), .CK(clk), .Q(
        pipeline_regfile_data[138]) );
  DFF_X1 pipeline_regfile_data_reg_5__10_ ( .D(n5253), .CK(clk), .Q(
        pipeline_regfile_data[170]) );
  DFF_X1 pipeline_regfile_data_reg_6__10_ ( .D(n5254), .CK(clk), .Q(
        pipeline_regfile_data[202]) );
  DFF_X1 pipeline_regfile_data_reg_7__10_ ( .D(n5255), .CK(clk), .Q(
        pipeline_regfile_data[234]) );
  DFF_X1 pipeline_regfile_data_reg_8__10_ ( .D(n5256), .CK(clk), .Q(
        pipeline_regfile_data[266]) );
  DFF_X1 pipeline_regfile_data_reg_9__10_ ( .D(n5257), .CK(clk), .Q(
        pipeline_regfile_data[298]) );
  DFF_X1 pipeline_regfile_data_reg_10__10_ ( .D(n5258), .CK(clk), .Q(
        pipeline_regfile_data[330]) );
  DFF_X1 pipeline_regfile_data_reg_11__10_ ( .D(n5259), .CK(clk), .Q(
        pipeline_regfile_data[362]) );
  DFF_X1 pipeline_regfile_data_reg_12__10_ ( .D(n5260), .CK(clk), .Q(
        pipeline_regfile_data[394]) );
  DFF_X1 pipeline_regfile_data_reg_13__10_ ( .D(n5261), .CK(clk), .Q(
        pipeline_regfile_data[426]) );
  DFF_X1 pipeline_regfile_data_reg_14__10_ ( .D(n5262), .CK(clk), .Q(
        pipeline_regfile_data[458]) );
  DFF_X1 pipeline_regfile_data_reg_15__10_ ( .D(n5263), .CK(clk), .Q(
        pipeline_regfile_data[490]) );
  DFF_X1 pipeline_regfile_data_reg_16__10_ ( .D(n5264), .CK(clk), .Q(
        pipeline_regfile_data[522]) );
  DFF_X1 pipeline_regfile_data_reg_17__10_ ( .D(n5265), .CK(clk), .Q(
        pipeline_regfile_data[554]) );
  DFF_X1 pipeline_regfile_data_reg_18__10_ ( .D(n5266), .CK(clk), .Q(
        pipeline_regfile_data[586]) );
  DFF_X1 pipeline_regfile_data_reg_19__10_ ( .D(n5267), .CK(clk), .Q(
        pipeline_regfile_data[618]) );
  DFF_X1 pipeline_regfile_data_reg_20__10_ ( .D(n5268), .CK(clk), .Q(
        pipeline_regfile_data[650]) );
  DFF_X1 pipeline_regfile_data_reg_21__10_ ( .D(n5269), .CK(clk), .Q(
        pipeline_regfile_data[682]) );
  DFF_X1 pipeline_regfile_data_reg_22__10_ ( .D(n5270), .CK(clk), .Q(
        pipeline_regfile_data[714]) );
  DFF_X1 pipeline_regfile_data_reg_23__10_ ( .D(n5271), .CK(clk), .Q(
        pipeline_regfile_data[746]) );
  DFF_X1 pipeline_regfile_data_reg_24__10_ ( .D(n5272), .CK(clk), .Q(
        pipeline_regfile_data[778]) );
  DFF_X1 pipeline_regfile_data_reg_25__10_ ( .D(n5273), .CK(clk), .Q(
        pipeline_regfile_data[810]) );
  DFF_X1 pipeline_regfile_data_reg_26__10_ ( .D(n5274), .CK(clk), .Q(
        pipeline_regfile_data[842]) );
  DFF_X1 pipeline_regfile_data_reg_27__10_ ( .D(n5275), .CK(clk), .Q(
        pipeline_regfile_data[874]) );
  DFF_X1 pipeline_regfile_data_reg_28__10_ ( .D(n5276), .CK(clk), .Q(
        pipeline_regfile_data[906]) );
  DFF_X1 pipeline_regfile_data_reg_29__10_ ( .D(n5277), .CK(clk), .Q(
        pipeline_regfile_data[938]) );
  DFF_X1 pipeline_regfile_data_reg_30__10_ ( .D(n5278), .CK(clk), .Q(
        pipeline_regfile_data[970]) );
  DFF_X1 pipeline_regfile_data_reg_31__10_ ( .D(n5279), .CK(clk), .Q(
        pipeline_regfile_data[1002]) );
  DFF_X1 pipeline_csr_mtime_full_reg_43_ ( .D(pipeline_csr_N2144), .CK(clk), 
        .Q(pipeline_csr_mtime_full[43]), .QN(n6907) );
  DFF_X1 pipeline_csr_mtime_full_reg_11_ ( .D(pipeline_csr_N2112), .CK(clk), 
        .Q(pipeline_csr_mtime_full[11]) );
  DFF_X1 pipeline_csr_time_full_reg_43_ ( .D(pipeline_csr_N1995), .CK(clk), 
        .Q(pipeline_csr_time_full[43]) );
  DFF_X1 pipeline_csr_time_full_reg_11_ ( .D(pipeline_csr_N1963), .CK(clk), 
        .Q(pipeline_csr_time_full[11]), .QN(n6893) );
  DFF_X1 pipeline_csr_cycle_full_reg_43_ ( .D(pipeline_csr_N1931), .CK(clk), 
        .Q(pipeline_csr_cycle_full[43]) );
  DFF_X1 pipeline_csr_cycle_full_reg_11_ ( .D(pipeline_csr_N1899), .CK(clk), 
        .Q(pipeline_csr_cycle_full[11]) );
  DFF_X1 pipeline_regfile_data_reg_1__11_ ( .D(n5218), .CK(clk), .Q(
        pipeline_regfile_data[43]) );
  DFF_X1 pipeline_regfile_data_reg_2__11_ ( .D(n5219), .CK(clk), .Q(
        pipeline_regfile_data[75]) );
  DFF_X1 pipeline_regfile_data_reg_3__11_ ( .D(n5220), .CK(clk), .Q(
        pipeline_regfile_data[107]) );
  DFF_X1 pipeline_regfile_data_reg_4__11_ ( .D(n5221), .CK(clk), .Q(
        pipeline_regfile_data[139]) );
  DFF_X1 pipeline_regfile_data_reg_5__11_ ( .D(n5222), .CK(clk), .Q(
        pipeline_regfile_data[171]) );
  DFF_X1 pipeline_regfile_data_reg_6__11_ ( .D(n5223), .CK(clk), .Q(
        pipeline_regfile_data[203]) );
  DFF_X1 pipeline_regfile_data_reg_7__11_ ( .D(n5224), .CK(clk), .Q(
        pipeline_regfile_data[235]) );
  DFF_X1 pipeline_regfile_data_reg_8__11_ ( .D(n5225), .CK(clk), .Q(
        pipeline_regfile_data[267]) );
  DFF_X1 pipeline_regfile_data_reg_9__11_ ( .D(n5226), .CK(clk), .Q(
        pipeline_regfile_data[299]) );
  DFF_X1 pipeline_regfile_data_reg_10__11_ ( .D(n5227), .CK(clk), .Q(
        pipeline_regfile_data[331]) );
  DFF_X1 pipeline_regfile_data_reg_11__11_ ( .D(n5228), .CK(clk), .Q(
        pipeline_regfile_data[363]) );
  DFF_X1 pipeline_regfile_data_reg_12__11_ ( .D(n5229), .CK(clk), .Q(
        pipeline_regfile_data[395]) );
  DFF_X1 pipeline_regfile_data_reg_13__11_ ( .D(n5230), .CK(clk), .Q(
        pipeline_regfile_data[427]) );
  DFF_X1 pipeline_regfile_data_reg_14__11_ ( .D(n5231), .CK(clk), .Q(
        pipeline_regfile_data[459]) );
  DFF_X1 pipeline_regfile_data_reg_15__11_ ( .D(n5232), .CK(clk), .Q(
        pipeline_regfile_data[491]) );
  DFF_X1 pipeline_regfile_data_reg_16__11_ ( .D(n5233), .CK(clk), .Q(
        pipeline_regfile_data[523]) );
  DFF_X1 pipeline_regfile_data_reg_17__11_ ( .D(n5234), .CK(clk), .Q(
        pipeline_regfile_data[555]) );
  DFF_X1 pipeline_regfile_data_reg_18__11_ ( .D(n5235), .CK(clk), .Q(
        pipeline_regfile_data[587]) );
  DFF_X1 pipeline_regfile_data_reg_19__11_ ( .D(n5236), .CK(clk), .Q(
        pipeline_regfile_data[619]) );
  DFF_X1 pipeline_regfile_data_reg_20__11_ ( .D(n5237), .CK(clk), .Q(
        pipeline_regfile_data[651]) );
  DFF_X1 pipeline_regfile_data_reg_21__11_ ( .D(n5238), .CK(clk), .Q(
        pipeline_regfile_data[683]) );
  DFF_X1 pipeline_regfile_data_reg_22__11_ ( .D(n5239), .CK(clk), .Q(
        pipeline_regfile_data[715]) );
  DFF_X1 pipeline_regfile_data_reg_23__11_ ( .D(n5240), .CK(clk), .Q(
        pipeline_regfile_data[747]) );
  DFF_X1 pipeline_regfile_data_reg_24__11_ ( .D(n5241), .CK(clk), .Q(
        pipeline_regfile_data[779]) );
  DFF_X1 pipeline_regfile_data_reg_25__11_ ( .D(n5242), .CK(clk), .Q(
        pipeline_regfile_data[811]) );
  DFF_X1 pipeline_regfile_data_reg_26__11_ ( .D(n5243), .CK(clk), .Q(
        pipeline_regfile_data[843]) );
  DFF_X1 pipeline_regfile_data_reg_27__11_ ( .D(n5244), .CK(clk), .Q(
        pipeline_regfile_data[875]) );
  DFF_X1 pipeline_regfile_data_reg_28__11_ ( .D(n5245), .CK(clk), .Q(
        pipeline_regfile_data[907]) );
  DFF_X1 pipeline_regfile_data_reg_29__11_ ( .D(n5246), .CK(clk), .Q(
        pipeline_regfile_data[939]) );
  DFF_X1 pipeline_regfile_data_reg_30__11_ ( .D(n5247), .CK(clk), .Q(
        pipeline_regfile_data[971]) );
  DFF_X1 pipeline_regfile_data_reg_31__11_ ( .D(n5248), .CK(clk), .Q(
        pipeline_regfile_data[1003]) );
  DFF_X1 pipeline_csr_mtime_full_reg_44_ ( .D(pipeline_csr_N2145), .CK(clk), 
        .Q(pipeline_csr_mtime_full[44]), .QN(n6906) );
  DFF_X1 pipeline_csr_mtime_full_reg_12_ ( .D(pipeline_csr_N2113), .CK(clk), 
        .Q(pipeline_csr_mtime_full[12]) );
  DFF_X1 pipeline_csr_time_full_reg_44_ ( .D(pipeline_csr_N1996), .CK(clk), 
        .Q(pipeline_csr_time_full[44]) );
  DFF_X1 pipeline_csr_time_full_reg_12_ ( .D(pipeline_csr_N1964), .CK(clk), 
        .Q(pipeline_csr_time_full[12]), .QN(n6883) );
  DFF_X1 pipeline_csr_cycle_full_reg_44_ ( .D(pipeline_csr_N1932), .CK(clk), 
        .Q(pipeline_csr_cycle_full[44]) );
  DFF_X1 pipeline_csr_cycle_full_reg_12_ ( .D(pipeline_csr_N1900), .CK(clk), 
        .Q(pipeline_csr_cycle_full[12]) );
  DFF_X1 pipeline_regfile_data_reg_1__12_ ( .D(n5187), .CK(clk), .Q(
        pipeline_regfile_data[44]) );
  DFF_X1 pipeline_regfile_data_reg_2__12_ ( .D(n5188), .CK(clk), .Q(
        pipeline_regfile_data[76]) );
  DFF_X1 pipeline_regfile_data_reg_3__12_ ( .D(n5189), .CK(clk), .Q(
        pipeline_regfile_data[108]) );
  DFF_X1 pipeline_regfile_data_reg_4__12_ ( .D(n5190), .CK(clk), .Q(
        pipeline_regfile_data[140]) );
  DFF_X1 pipeline_regfile_data_reg_5__12_ ( .D(n5191), .CK(clk), .Q(
        pipeline_regfile_data[172]) );
  DFF_X1 pipeline_regfile_data_reg_6__12_ ( .D(n5192), .CK(clk), .Q(
        pipeline_regfile_data[204]) );
  DFF_X1 pipeline_regfile_data_reg_7__12_ ( .D(n5193), .CK(clk), .Q(
        pipeline_regfile_data[236]) );
  DFF_X1 pipeline_regfile_data_reg_8__12_ ( .D(n5194), .CK(clk), .Q(
        pipeline_regfile_data[268]) );
  DFF_X1 pipeline_regfile_data_reg_9__12_ ( .D(n5195), .CK(clk), .Q(
        pipeline_regfile_data[300]) );
  DFF_X1 pipeline_regfile_data_reg_10__12_ ( .D(n5196), .CK(clk), .Q(
        pipeline_regfile_data[332]) );
  DFF_X1 pipeline_regfile_data_reg_11__12_ ( .D(n5197), .CK(clk), .Q(
        pipeline_regfile_data[364]) );
  DFF_X1 pipeline_regfile_data_reg_12__12_ ( .D(n5198), .CK(clk), .Q(
        pipeline_regfile_data[396]) );
  DFF_X1 pipeline_regfile_data_reg_13__12_ ( .D(n5199), .CK(clk), .Q(
        pipeline_regfile_data[428]) );
  DFF_X1 pipeline_regfile_data_reg_14__12_ ( .D(n5200), .CK(clk), .Q(
        pipeline_regfile_data[460]) );
  DFF_X1 pipeline_regfile_data_reg_15__12_ ( .D(n5201), .CK(clk), .Q(
        pipeline_regfile_data[492]) );
  DFF_X1 pipeline_regfile_data_reg_16__12_ ( .D(n5202), .CK(clk), .Q(
        pipeline_regfile_data[524]) );
  DFF_X1 pipeline_regfile_data_reg_17__12_ ( .D(n5203), .CK(clk), .Q(
        pipeline_regfile_data[556]) );
  DFF_X1 pipeline_regfile_data_reg_18__12_ ( .D(n5204), .CK(clk), .Q(
        pipeline_regfile_data[588]) );
  DFF_X1 pipeline_regfile_data_reg_19__12_ ( .D(n5205), .CK(clk), .Q(
        pipeline_regfile_data[620]) );
  DFF_X1 pipeline_regfile_data_reg_20__12_ ( .D(n5206), .CK(clk), .Q(
        pipeline_regfile_data[652]) );
  DFF_X1 pipeline_regfile_data_reg_21__12_ ( .D(n5207), .CK(clk), .Q(
        pipeline_regfile_data[684]) );
  DFF_X1 pipeline_regfile_data_reg_22__12_ ( .D(n5208), .CK(clk), .Q(
        pipeline_regfile_data[716]) );
  DFF_X1 pipeline_regfile_data_reg_23__12_ ( .D(n5209), .CK(clk), .Q(
        pipeline_regfile_data[748]) );
  DFF_X1 pipeline_regfile_data_reg_24__12_ ( .D(n5210), .CK(clk), .Q(
        pipeline_regfile_data[780]) );
  DFF_X1 pipeline_regfile_data_reg_25__12_ ( .D(n5211), .CK(clk), .Q(
        pipeline_regfile_data[812]) );
  DFF_X1 pipeline_regfile_data_reg_26__12_ ( .D(n5212), .CK(clk), .Q(
        pipeline_regfile_data[844]) );
  DFF_X1 pipeline_regfile_data_reg_27__12_ ( .D(n5213), .CK(clk), .Q(
        pipeline_regfile_data[876]) );
  DFF_X1 pipeline_regfile_data_reg_28__12_ ( .D(n5214), .CK(clk), .Q(
        pipeline_regfile_data[908]) );
  DFF_X1 pipeline_regfile_data_reg_29__12_ ( .D(n5215), .CK(clk), .Q(
        pipeline_regfile_data[940]) );
  DFF_X1 pipeline_regfile_data_reg_30__12_ ( .D(n5216), .CK(clk), .Q(
        pipeline_regfile_data[972]) );
  DFF_X1 pipeline_regfile_data_reg_31__12_ ( .D(n5217), .CK(clk), .Q(
        pipeline_regfile_data[1004]) );
  DFF_X1 pipeline_csr_mtime_full_reg_45_ ( .D(pipeline_csr_N2146), .CK(clk), 
        .Q(pipeline_csr_mtime_full[45]), .QN(n6905) );
  DFF_X1 pipeline_csr_mtime_full_reg_13_ ( .D(pipeline_csr_N2114), .CK(clk), 
        .Q(pipeline_csr_mtime_full[13]) );
  DFF_X1 pipeline_csr_time_full_reg_45_ ( .D(pipeline_csr_N1997), .CK(clk), 
        .Q(pipeline_csr_time_full[45]) );
  DFF_X1 pipeline_csr_time_full_reg_13_ ( .D(pipeline_csr_N1965), .CK(clk), 
        .Q(pipeline_csr_time_full[13]), .QN(n6895) );
  DFF_X1 pipeline_csr_cycle_full_reg_45_ ( .D(pipeline_csr_N1933), .CK(clk), 
        .Q(pipeline_csr_cycle_full[45]) );
  DFF_X1 pipeline_csr_cycle_full_reg_13_ ( .D(pipeline_csr_N1901), .CK(clk), 
        .Q(pipeline_csr_cycle_full[13]) );
  DFF_X1 pipeline_regfile_data_reg_1__13_ ( .D(n5156), .CK(clk), .Q(
        pipeline_regfile_data[45]) );
  DFF_X1 pipeline_regfile_data_reg_2__13_ ( .D(n5157), .CK(clk), .Q(
        pipeline_regfile_data[77]) );
  DFF_X1 pipeline_regfile_data_reg_3__13_ ( .D(n5158), .CK(clk), .Q(
        pipeline_regfile_data[109]) );
  DFF_X1 pipeline_regfile_data_reg_4__13_ ( .D(n5159), .CK(clk), .Q(
        pipeline_regfile_data[141]) );
  DFF_X1 pipeline_regfile_data_reg_5__13_ ( .D(n5160), .CK(clk), .Q(
        pipeline_regfile_data[173]) );
  DFF_X1 pipeline_regfile_data_reg_6__13_ ( .D(n5161), .CK(clk), .Q(
        pipeline_regfile_data[205]) );
  DFF_X1 pipeline_regfile_data_reg_7__13_ ( .D(n5162), .CK(clk), .Q(
        pipeline_regfile_data[237]) );
  DFF_X1 pipeline_regfile_data_reg_8__13_ ( .D(n5163), .CK(clk), .Q(
        pipeline_regfile_data[269]) );
  DFF_X1 pipeline_regfile_data_reg_9__13_ ( .D(n5164), .CK(clk), .Q(
        pipeline_regfile_data[301]) );
  DFF_X1 pipeline_regfile_data_reg_10__13_ ( .D(n5165), .CK(clk), .Q(
        pipeline_regfile_data[333]) );
  DFF_X1 pipeline_regfile_data_reg_11__13_ ( .D(n5166), .CK(clk), .Q(
        pipeline_regfile_data[365]) );
  DFF_X1 pipeline_regfile_data_reg_12__13_ ( .D(n5167), .CK(clk), .Q(
        pipeline_regfile_data[397]) );
  DFF_X1 pipeline_regfile_data_reg_13__13_ ( .D(n5168), .CK(clk), .Q(
        pipeline_regfile_data[429]) );
  DFF_X1 pipeline_regfile_data_reg_14__13_ ( .D(n5169), .CK(clk), .Q(
        pipeline_regfile_data[461]) );
  DFF_X1 pipeline_regfile_data_reg_15__13_ ( .D(n5170), .CK(clk), .Q(
        pipeline_regfile_data[493]) );
  DFF_X1 pipeline_regfile_data_reg_16__13_ ( .D(n5171), .CK(clk), .Q(
        pipeline_regfile_data[525]) );
  DFF_X1 pipeline_regfile_data_reg_17__13_ ( .D(n5172), .CK(clk), .Q(
        pipeline_regfile_data[557]) );
  DFF_X1 pipeline_regfile_data_reg_18__13_ ( .D(n5173), .CK(clk), .Q(
        pipeline_regfile_data[589]) );
  DFF_X1 pipeline_regfile_data_reg_19__13_ ( .D(n5174), .CK(clk), .Q(
        pipeline_regfile_data[621]) );
  DFF_X1 pipeline_regfile_data_reg_20__13_ ( .D(n5175), .CK(clk), .Q(
        pipeline_regfile_data[653]) );
  DFF_X1 pipeline_regfile_data_reg_21__13_ ( .D(n5176), .CK(clk), .Q(
        pipeline_regfile_data[685]) );
  DFF_X1 pipeline_regfile_data_reg_22__13_ ( .D(n5177), .CK(clk), .Q(
        pipeline_regfile_data[717]) );
  DFF_X1 pipeline_regfile_data_reg_23__13_ ( .D(n5178), .CK(clk), .Q(
        pipeline_regfile_data[749]) );
  DFF_X1 pipeline_regfile_data_reg_24__13_ ( .D(n5179), .CK(clk), .Q(
        pipeline_regfile_data[781]) );
  DFF_X1 pipeline_regfile_data_reg_25__13_ ( .D(n5180), .CK(clk), .Q(
        pipeline_regfile_data[813]) );
  DFF_X1 pipeline_regfile_data_reg_26__13_ ( .D(n5181), .CK(clk), .Q(
        pipeline_regfile_data[845]) );
  DFF_X1 pipeline_regfile_data_reg_27__13_ ( .D(n5182), .CK(clk), .Q(
        pipeline_regfile_data[877]) );
  DFF_X1 pipeline_regfile_data_reg_28__13_ ( .D(n5183), .CK(clk), .Q(
        pipeline_regfile_data[909]) );
  DFF_X1 pipeline_regfile_data_reg_29__13_ ( .D(n5184), .CK(clk), .Q(
        pipeline_regfile_data[941]) );
  DFF_X1 pipeline_regfile_data_reg_30__13_ ( .D(n5185), .CK(clk), .Q(
        pipeline_regfile_data[973]) );
  DFF_X1 pipeline_regfile_data_reg_31__13_ ( .D(n5186), .CK(clk), .Q(
        pipeline_regfile_data[1005]) );
  DFF_X1 pipeline_csr_mtime_full_reg_46_ ( .D(pipeline_csr_N2147), .CK(clk), 
        .Q(pipeline_csr_mtime_full[46]), .QN(n6904) );
  DFF_X1 pipeline_csr_mtime_full_reg_14_ ( .D(pipeline_csr_N2115), .CK(clk), 
        .Q(pipeline_csr_mtime_full[14]), .QN(n6858) );
  DFF_X1 pipeline_csr_time_full_reg_46_ ( .D(pipeline_csr_N1998), .CK(clk), 
        .Q(pipeline_csr_time_full[46]) );
  DFF_X1 pipeline_csr_time_full_reg_14_ ( .D(pipeline_csr_N1966), .CK(clk), 
        .Q(pipeline_csr_time_full[14]), .QN(n6886) );
  DFF_X1 pipeline_csr_cycle_full_reg_46_ ( .D(pipeline_csr_N1934), .CK(clk), 
        .Q(pipeline_csr_cycle_full[46]) );
  DFF_X1 pipeline_csr_cycle_full_reg_14_ ( .D(pipeline_csr_N1902), .CK(clk), 
        .Q(pipeline_csr_cycle_full[14]) );
  DFF_X1 pipeline_regfile_data_reg_1__14_ ( .D(n5125), .CK(clk), .Q(
        pipeline_regfile_data[46]) );
  DFF_X1 pipeline_regfile_data_reg_2__14_ ( .D(n5126), .CK(clk), .Q(
        pipeline_regfile_data[78]) );
  DFF_X1 pipeline_regfile_data_reg_3__14_ ( .D(n5127), .CK(clk), .Q(
        pipeline_regfile_data[110]) );
  DFF_X1 pipeline_regfile_data_reg_4__14_ ( .D(n5128), .CK(clk), .Q(
        pipeline_regfile_data[142]) );
  DFF_X1 pipeline_regfile_data_reg_5__14_ ( .D(n5129), .CK(clk), .Q(
        pipeline_regfile_data[174]) );
  DFF_X1 pipeline_regfile_data_reg_6__14_ ( .D(n5130), .CK(clk), .Q(
        pipeline_regfile_data[206]) );
  DFF_X1 pipeline_regfile_data_reg_7__14_ ( .D(n5131), .CK(clk), .Q(
        pipeline_regfile_data[238]) );
  DFF_X1 pipeline_regfile_data_reg_8__14_ ( .D(n5132), .CK(clk), .Q(
        pipeline_regfile_data[270]) );
  DFF_X1 pipeline_regfile_data_reg_9__14_ ( .D(n5133), .CK(clk), .Q(
        pipeline_regfile_data[302]) );
  DFF_X1 pipeline_regfile_data_reg_10__14_ ( .D(n5134), .CK(clk), .Q(
        pipeline_regfile_data[334]) );
  DFF_X1 pipeline_regfile_data_reg_11__14_ ( .D(n5135), .CK(clk), .Q(
        pipeline_regfile_data[366]) );
  DFF_X1 pipeline_regfile_data_reg_12__14_ ( .D(n5136), .CK(clk), .Q(
        pipeline_regfile_data[398]) );
  DFF_X1 pipeline_regfile_data_reg_13__14_ ( .D(n5137), .CK(clk), .Q(
        pipeline_regfile_data[430]) );
  DFF_X1 pipeline_regfile_data_reg_14__14_ ( .D(n5138), .CK(clk), .Q(
        pipeline_regfile_data[462]) );
  DFF_X1 pipeline_regfile_data_reg_15__14_ ( .D(n5139), .CK(clk), .Q(
        pipeline_regfile_data[494]) );
  DFF_X1 pipeline_regfile_data_reg_16__14_ ( .D(n5140), .CK(clk), .Q(
        pipeline_regfile_data[526]) );
  DFF_X1 pipeline_regfile_data_reg_17__14_ ( .D(n5141), .CK(clk), .Q(
        pipeline_regfile_data[558]) );
  DFF_X1 pipeline_regfile_data_reg_18__14_ ( .D(n5142), .CK(clk), .Q(
        pipeline_regfile_data[590]) );
  DFF_X1 pipeline_regfile_data_reg_19__14_ ( .D(n5143), .CK(clk), .Q(
        pipeline_regfile_data[622]) );
  DFF_X1 pipeline_regfile_data_reg_20__14_ ( .D(n5144), .CK(clk), .Q(
        pipeline_regfile_data[654]) );
  DFF_X1 pipeline_regfile_data_reg_21__14_ ( .D(n5145), .CK(clk), .Q(
        pipeline_regfile_data[686]) );
  DFF_X1 pipeline_regfile_data_reg_22__14_ ( .D(n5146), .CK(clk), .Q(
        pipeline_regfile_data[718]) );
  DFF_X1 pipeline_regfile_data_reg_23__14_ ( .D(n5147), .CK(clk), .Q(
        pipeline_regfile_data[750]) );
  DFF_X1 pipeline_regfile_data_reg_24__14_ ( .D(n5148), .CK(clk), .Q(
        pipeline_regfile_data[782]) );
  DFF_X1 pipeline_regfile_data_reg_25__14_ ( .D(n5149), .CK(clk), .Q(
        pipeline_regfile_data[814]) );
  DFF_X1 pipeline_regfile_data_reg_26__14_ ( .D(n5150), .CK(clk), .Q(
        pipeline_regfile_data[846]) );
  DFF_X1 pipeline_regfile_data_reg_27__14_ ( .D(n5151), .CK(clk), .Q(
        pipeline_regfile_data[878]) );
  DFF_X1 pipeline_regfile_data_reg_28__14_ ( .D(n5152), .CK(clk), .Q(
        pipeline_regfile_data[910]) );
  DFF_X1 pipeline_regfile_data_reg_29__14_ ( .D(n5153), .CK(clk), .Q(
        pipeline_regfile_data[942]) );
  DFF_X1 pipeline_regfile_data_reg_30__14_ ( .D(n5154), .CK(clk), .Q(
        pipeline_regfile_data[974]) );
  DFF_X1 pipeline_regfile_data_reg_31__14_ ( .D(n5155), .CK(clk), .Q(
        pipeline_regfile_data[1006]) );
  DFF_X1 pipeline_csr_mtime_full_reg_47_ ( .D(pipeline_csr_N2148), .CK(clk), 
        .Q(pipeline_csr_mtime_full[47]) );
  DFF_X2 pipeline_csr_instret_full_reg_47_ ( .D(n5999), .CK(clk), .Q(n11104), 
        .QN(n1430) );
  DFF_X1 pipeline_csr_mtime_full_reg_15_ ( .D(pipeline_csr_N2116), .CK(clk), 
        .Q(pipeline_csr_mtime_full[15]), .QN(n6865) );
  DFF_X1 pipeline_csr_time_full_reg_15_ ( .D(pipeline_csr_N1967), .CK(clk), 
        .Q(pipeline_csr_time_full[15]) );
  DFF_X1 pipeline_csr_cycle_full_reg_47_ ( .D(pipeline_csr_N1935), .CK(clk), 
        .Q(pipeline_csr_cycle_full[47]), .QN(n6882) );
  DFF_X1 pipeline_csr_cycle_full_reg_15_ ( .D(pipeline_csr_N1903), .CK(clk), 
        .Q(pipeline_csr_cycle_full[15]) );
  DFF_X1 pipeline_regfile_data_reg_1__15_ ( .D(n5094), .CK(clk), .Q(
        pipeline_regfile_data[47]) );
  DFF_X1 pipeline_regfile_data_reg_2__15_ ( .D(n5095), .CK(clk), .Q(
        pipeline_regfile_data[79]) );
  DFF_X1 pipeline_regfile_data_reg_3__15_ ( .D(n5096), .CK(clk), .Q(
        pipeline_regfile_data[111]) );
  DFF_X1 pipeline_regfile_data_reg_4__15_ ( .D(n5097), .CK(clk), .Q(
        pipeline_regfile_data[143]) );
  DFF_X1 pipeline_regfile_data_reg_5__15_ ( .D(n5098), .CK(clk), .Q(
        pipeline_regfile_data[175]) );
  DFF_X1 pipeline_regfile_data_reg_6__15_ ( .D(n5099), .CK(clk), .Q(
        pipeline_regfile_data[207]) );
  DFF_X1 pipeline_regfile_data_reg_7__15_ ( .D(n5100), .CK(clk), .Q(
        pipeline_regfile_data[239]) );
  DFF_X1 pipeline_regfile_data_reg_8__15_ ( .D(n5101), .CK(clk), .Q(
        pipeline_regfile_data[271]) );
  DFF_X1 pipeline_regfile_data_reg_9__15_ ( .D(n5102), .CK(clk), .Q(
        pipeline_regfile_data[303]) );
  DFF_X1 pipeline_regfile_data_reg_10__15_ ( .D(n5103), .CK(clk), .Q(
        pipeline_regfile_data[335]) );
  DFF_X1 pipeline_regfile_data_reg_11__15_ ( .D(n5104), .CK(clk), .Q(
        pipeline_regfile_data[367]) );
  DFF_X1 pipeline_regfile_data_reg_12__15_ ( .D(n5105), .CK(clk), .Q(
        pipeline_regfile_data[399]) );
  DFF_X1 pipeline_regfile_data_reg_13__15_ ( .D(n5106), .CK(clk), .Q(
        pipeline_regfile_data[431]) );
  DFF_X1 pipeline_regfile_data_reg_14__15_ ( .D(n5107), .CK(clk), .Q(
        pipeline_regfile_data[463]) );
  DFF_X1 pipeline_regfile_data_reg_15__15_ ( .D(n5108), .CK(clk), .Q(
        pipeline_regfile_data[495]) );
  DFF_X1 pipeline_regfile_data_reg_16__15_ ( .D(n5109), .CK(clk), .Q(
        pipeline_regfile_data[527]) );
  DFF_X1 pipeline_regfile_data_reg_17__15_ ( .D(n5110), .CK(clk), .Q(
        pipeline_regfile_data[559]) );
  DFF_X1 pipeline_regfile_data_reg_18__15_ ( .D(n5111), .CK(clk), .Q(
        pipeline_regfile_data[591]) );
  DFF_X1 pipeline_regfile_data_reg_19__15_ ( .D(n5112), .CK(clk), .Q(
        pipeline_regfile_data[623]) );
  DFF_X1 pipeline_regfile_data_reg_20__15_ ( .D(n5113), .CK(clk), .Q(
        pipeline_regfile_data[655]) );
  DFF_X1 pipeline_regfile_data_reg_21__15_ ( .D(n5114), .CK(clk), .Q(
        pipeline_regfile_data[687]) );
  DFF_X1 pipeline_regfile_data_reg_22__15_ ( .D(n5115), .CK(clk), .Q(
        pipeline_regfile_data[719]) );
  DFF_X1 pipeline_regfile_data_reg_23__15_ ( .D(n5116), .CK(clk), .Q(
        pipeline_regfile_data[751]) );
  DFF_X1 pipeline_regfile_data_reg_24__15_ ( .D(n5117), .CK(clk), .Q(
        pipeline_regfile_data[783]) );
  DFF_X1 pipeline_regfile_data_reg_25__15_ ( .D(n5118), .CK(clk), .Q(
        pipeline_regfile_data[815]) );
  DFF_X1 pipeline_regfile_data_reg_26__15_ ( .D(n5119), .CK(clk), .Q(
        pipeline_regfile_data[847]) );
  DFF_X1 pipeline_regfile_data_reg_27__15_ ( .D(n5120), .CK(clk), .Q(
        pipeline_regfile_data[879]) );
  DFF_X1 pipeline_regfile_data_reg_28__15_ ( .D(n5121), .CK(clk), .Q(
        pipeline_regfile_data[911]) );
  DFF_X1 pipeline_regfile_data_reg_29__15_ ( .D(n5122), .CK(clk), .Q(
        pipeline_regfile_data[943]) );
  DFF_X1 pipeline_regfile_data_reg_30__15_ ( .D(n5123), .CK(clk), .Q(
        pipeline_regfile_data[975]) );
  DFF_X1 pipeline_regfile_data_reg_31__15_ ( .D(n5124), .CK(clk), .Q(
        pipeline_regfile_data[1007]) );
  DFF_X1 pipeline_csr_mtime_full_reg_48_ ( .D(pipeline_csr_N2149), .CK(clk), 
        .Q(pipeline_csr_mtime_full[48]), .QN(n6903) );
  DFF_X1 pipeline_csr_mtime_full_reg_16_ ( .D(pipeline_csr_N2117), .CK(clk), 
        .Q(pipeline_csr_mtime_full[16]), .QN(n6857) );
  DFF_X1 pipeline_csr_time_full_reg_48_ ( .D(pipeline_csr_N2000), .CK(clk), 
        .Q(pipeline_csr_time_full[48]) );
  DFF_X1 pipeline_csr_time_full_reg_16_ ( .D(pipeline_csr_N1968), .CK(clk), 
        .Q(pipeline_csr_time_full[16]), .QN(n6885) );
  DFF_X1 pipeline_csr_cycle_full_reg_48_ ( .D(pipeline_csr_N1936), .CK(clk), 
        .Q(pipeline_csr_cycle_full[48]) );
  DFF_X1 pipeline_csr_cycle_full_reg_16_ ( .D(pipeline_csr_N1904), .CK(clk), 
        .Q(pipeline_csr_cycle_full[16]) );
  DFF_X1 pipeline_regfile_data_reg_1__16_ ( .D(n5063), .CK(clk), .Q(
        pipeline_regfile_data[48]) );
  DFF_X1 pipeline_regfile_data_reg_2__16_ ( .D(n5064), .CK(clk), .Q(
        pipeline_regfile_data[80]) );
  DFF_X1 pipeline_regfile_data_reg_3__16_ ( .D(n5065), .CK(clk), .Q(
        pipeline_regfile_data[112]) );
  DFF_X1 pipeline_regfile_data_reg_4__16_ ( .D(n5066), .CK(clk), .Q(
        pipeline_regfile_data[144]) );
  DFF_X1 pipeline_regfile_data_reg_5__16_ ( .D(n5067), .CK(clk), .Q(
        pipeline_regfile_data[176]) );
  DFF_X1 pipeline_regfile_data_reg_6__16_ ( .D(n5068), .CK(clk), .Q(
        pipeline_regfile_data[208]) );
  DFF_X1 pipeline_regfile_data_reg_7__16_ ( .D(n5069), .CK(clk), .Q(
        pipeline_regfile_data[240]) );
  DFF_X1 pipeline_regfile_data_reg_8__16_ ( .D(n5070), .CK(clk), .Q(
        pipeline_regfile_data[272]) );
  DFF_X1 pipeline_regfile_data_reg_9__16_ ( .D(n5071), .CK(clk), .Q(
        pipeline_regfile_data[304]) );
  DFF_X1 pipeline_regfile_data_reg_10__16_ ( .D(n5072), .CK(clk), .Q(
        pipeline_regfile_data[336]) );
  DFF_X1 pipeline_regfile_data_reg_11__16_ ( .D(n5073), .CK(clk), .Q(
        pipeline_regfile_data[368]) );
  DFF_X1 pipeline_regfile_data_reg_12__16_ ( .D(n5074), .CK(clk), .Q(
        pipeline_regfile_data[400]) );
  DFF_X1 pipeline_regfile_data_reg_13__16_ ( .D(n5075), .CK(clk), .Q(
        pipeline_regfile_data[432]) );
  DFF_X1 pipeline_regfile_data_reg_14__16_ ( .D(n5076), .CK(clk), .Q(
        pipeline_regfile_data[464]) );
  DFF_X1 pipeline_regfile_data_reg_15__16_ ( .D(n5077), .CK(clk), .Q(
        pipeline_regfile_data[496]) );
  DFF_X1 pipeline_regfile_data_reg_16__16_ ( .D(n5078), .CK(clk), .Q(
        pipeline_regfile_data[528]) );
  DFF_X1 pipeline_regfile_data_reg_17__16_ ( .D(n5079), .CK(clk), .Q(
        pipeline_regfile_data[560]) );
  DFF_X1 pipeline_regfile_data_reg_18__16_ ( .D(n5080), .CK(clk), .Q(
        pipeline_regfile_data[592]) );
  DFF_X1 pipeline_regfile_data_reg_19__16_ ( .D(n5081), .CK(clk), .Q(
        pipeline_regfile_data[624]) );
  DFF_X1 pipeline_regfile_data_reg_20__16_ ( .D(n5082), .CK(clk), .Q(
        pipeline_regfile_data[656]) );
  DFF_X1 pipeline_regfile_data_reg_21__16_ ( .D(n5083), .CK(clk), .Q(
        pipeline_regfile_data[688]) );
  DFF_X1 pipeline_regfile_data_reg_22__16_ ( .D(n5084), .CK(clk), .Q(
        pipeline_regfile_data[720]) );
  DFF_X1 pipeline_regfile_data_reg_23__16_ ( .D(n5085), .CK(clk), .Q(
        pipeline_regfile_data[752]) );
  DFF_X1 pipeline_regfile_data_reg_24__16_ ( .D(n5086), .CK(clk), .Q(
        pipeline_regfile_data[784]) );
  DFF_X1 pipeline_regfile_data_reg_25__16_ ( .D(n5087), .CK(clk), .Q(
        pipeline_regfile_data[816]) );
  DFF_X1 pipeline_regfile_data_reg_26__16_ ( .D(n5088), .CK(clk), .Q(
        pipeline_regfile_data[848]) );
  DFF_X1 pipeline_regfile_data_reg_27__16_ ( .D(n5089), .CK(clk), .Q(
        pipeline_regfile_data[880]) );
  DFF_X1 pipeline_regfile_data_reg_28__16_ ( .D(n5090), .CK(clk), .Q(
        pipeline_regfile_data[912]) );
  DFF_X1 pipeline_regfile_data_reg_29__16_ ( .D(n5091), .CK(clk), .Q(
        pipeline_regfile_data[944]) );
  DFF_X1 pipeline_regfile_data_reg_30__16_ ( .D(n5092), .CK(clk), .Q(
        pipeline_regfile_data[976]) );
  DFF_X1 pipeline_regfile_data_reg_31__16_ ( .D(n5093), .CK(clk), .Q(
        pipeline_regfile_data[1008]) );
  DFF_X1 pipeline_csr_mtime_full_reg_49_ ( .D(pipeline_csr_N2150), .CK(clk), 
        .Q(pipeline_csr_mtime_full[49]), .QN(n6902) );
  DFF_X1 pipeline_csr_mtime_full_reg_17_ ( .D(pipeline_csr_N2118), .CK(clk), 
        .Q(pipeline_csr_mtime_full[17]) );
  DFF_X1 pipeline_csr_time_full_reg_49_ ( .D(pipeline_csr_N2001), .CK(clk), 
        .Q(pipeline_csr_time_full[49]) );
  DFF_X1 pipeline_csr_time_full_reg_17_ ( .D(pipeline_csr_N1969), .CK(clk), 
        .Q(pipeline_csr_time_full[17]), .QN(n6896) );
  DFF_X1 pipeline_csr_cycle_full_reg_49_ ( .D(pipeline_csr_N1937), .CK(clk), 
        .Q(pipeline_csr_cycle_full[49]) );
  DFF_X1 pipeline_csr_cycle_full_reg_17_ ( .D(pipeline_csr_N1905), .CK(clk), 
        .Q(pipeline_csr_cycle_full[17]) );
  DFF_X1 pipeline_regfile_data_reg_1__17_ ( .D(n5032), .CK(clk), .Q(
        pipeline_regfile_data[49]) );
  DFF_X1 pipeline_regfile_data_reg_2__17_ ( .D(n5033), .CK(clk), .Q(
        pipeline_regfile_data[81]) );
  DFF_X1 pipeline_regfile_data_reg_3__17_ ( .D(n5034), .CK(clk), .Q(
        pipeline_regfile_data[113]) );
  DFF_X1 pipeline_regfile_data_reg_4__17_ ( .D(n5035), .CK(clk), .Q(
        pipeline_regfile_data[145]) );
  DFF_X1 pipeline_regfile_data_reg_5__17_ ( .D(n5036), .CK(clk), .Q(
        pipeline_regfile_data[177]) );
  DFF_X1 pipeline_regfile_data_reg_6__17_ ( .D(n5037), .CK(clk), .Q(
        pipeline_regfile_data[209]) );
  DFF_X1 pipeline_regfile_data_reg_7__17_ ( .D(n5038), .CK(clk), .Q(
        pipeline_regfile_data[241]) );
  DFF_X1 pipeline_regfile_data_reg_8__17_ ( .D(n5039), .CK(clk), .Q(
        pipeline_regfile_data[273]) );
  DFF_X1 pipeline_regfile_data_reg_9__17_ ( .D(n5040), .CK(clk), .Q(
        pipeline_regfile_data[305]) );
  DFF_X1 pipeline_regfile_data_reg_10__17_ ( .D(n5041), .CK(clk), .Q(
        pipeline_regfile_data[337]) );
  DFF_X1 pipeline_regfile_data_reg_11__17_ ( .D(n5042), .CK(clk), .Q(
        pipeline_regfile_data[369]) );
  DFF_X1 pipeline_regfile_data_reg_12__17_ ( .D(n5043), .CK(clk), .Q(
        pipeline_regfile_data[401]) );
  DFF_X1 pipeline_regfile_data_reg_13__17_ ( .D(n5044), .CK(clk), .Q(
        pipeline_regfile_data[433]) );
  DFF_X1 pipeline_regfile_data_reg_14__17_ ( .D(n5045), .CK(clk), .Q(
        pipeline_regfile_data[465]) );
  DFF_X1 pipeline_regfile_data_reg_15__17_ ( .D(n5046), .CK(clk), .Q(
        pipeline_regfile_data[497]) );
  DFF_X1 pipeline_regfile_data_reg_16__17_ ( .D(n5047), .CK(clk), .Q(
        pipeline_regfile_data[529]) );
  DFF_X1 pipeline_regfile_data_reg_17__17_ ( .D(n5048), .CK(clk), .Q(
        pipeline_regfile_data[561]) );
  DFF_X1 pipeline_regfile_data_reg_18__17_ ( .D(n5049), .CK(clk), .Q(
        pipeline_regfile_data[593]) );
  DFF_X1 pipeline_regfile_data_reg_19__17_ ( .D(n5050), .CK(clk), .Q(
        pipeline_regfile_data[625]) );
  DFF_X1 pipeline_regfile_data_reg_20__17_ ( .D(n5051), .CK(clk), .Q(
        pipeline_regfile_data[657]) );
  DFF_X1 pipeline_regfile_data_reg_21__17_ ( .D(n5052), .CK(clk), .Q(
        pipeline_regfile_data[689]) );
  DFF_X1 pipeline_regfile_data_reg_22__17_ ( .D(n5053), .CK(clk), .Q(
        pipeline_regfile_data[721]) );
  DFF_X1 pipeline_regfile_data_reg_23__17_ ( .D(n5054), .CK(clk), .Q(
        pipeline_regfile_data[753]) );
  DFF_X1 pipeline_regfile_data_reg_24__17_ ( .D(n5055), .CK(clk), .Q(
        pipeline_regfile_data[785]) );
  DFF_X1 pipeline_regfile_data_reg_25__17_ ( .D(n5056), .CK(clk), .Q(
        pipeline_regfile_data[817]) );
  DFF_X1 pipeline_regfile_data_reg_26__17_ ( .D(n5057), .CK(clk), .Q(
        pipeline_regfile_data[849]) );
  DFF_X1 pipeline_regfile_data_reg_27__17_ ( .D(n5058), .CK(clk), .Q(
        pipeline_regfile_data[881]) );
  DFF_X1 pipeline_regfile_data_reg_28__17_ ( .D(n5059), .CK(clk), .Q(
        pipeline_regfile_data[913]) );
  DFF_X1 pipeline_regfile_data_reg_29__17_ ( .D(n5060), .CK(clk), .Q(
        pipeline_regfile_data[945]) );
  DFF_X1 pipeline_regfile_data_reg_30__17_ ( .D(n5061), .CK(clk), .Q(
        pipeline_regfile_data[977]) );
  DFF_X1 pipeline_regfile_data_reg_31__17_ ( .D(n5062), .CK(clk), .Q(
        pipeline_regfile_data[1009]) );
  DFF_X1 pipeline_csr_mtime_full_reg_50_ ( .D(pipeline_csr_N2151), .CK(clk), 
        .Q(pipeline_csr_mtime_full[50]), .QN(n6881) );
  DFF_X1 pipeline_csr_mtime_full_reg_18_ ( .D(pipeline_csr_N2119), .CK(clk), 
        .Q(pipeline_csr_mtime_full[18]), .QN(n6851) );
  DFF_X1 pipeline_csr_time_full_reg_50_ ( .D(pipeline_csr_N2002), .CK(clk), 
        .Q(pipeline_csr_time_full[50]) );
  DFF_X1 pipeline_csr_time_full_reg_18_ ( .D(pipeline_csr_N1970), .CK(clk), 
        .Q(pipeline_csr_time_full[18]), .QN(n6864) );
  DFF_X1 pipeline_csr_cycle_full_reg_50_ ( .D(pipeline_csr_N1938), .CK(clk), 
        .Q(pipeline_csr_cycle_full[50]) );
  DFF_X1 pipeline_csr_cycle_full_reg_18_ ( .D(pipeline_csr_N1906), .CK(clk), 
        .Q(pipeline_csr_cycle_full[18]) );
  DFF_X1 pipeline_regfile_data_reg_1__18_ ( .D(n5001), .CK(clk), .Q(
        pipeline_regfile_data[50]) );
  DFF_X1 pipeline_regfile_data_reg_2__18_ ( .D(n5002), .CK(clk), .Q(
        pipeline_regfile_data[82]) );
  DFF_X1 pipeline_regfile_data_reg_3__18_ ( .D(n5003), .CK(clk), .Q(
        pipeline_regfile_data[114]) );
  DFF_X1 pipeline_regfile_data_reg_4__18_ ( .D(n5004), .CK(clk), .Q(
        pipeline_regfile_data[146]) );
  DFF_X1 pipeline_regfile_data_reg_5__18_ ( .D(n5005), .CK(clk), .Q(
        pipeline_regfile_data[178]) );
  DFF_X1 pipeline_regfile_data_reg_6__18_ ( .D(n5006), .CK(clk), .Q(
        pipeline_regfile_data[210]) );
  DFF_X1 pipeline_regfile_data_reg_7__18_ ( .D(n5007), .CK(clk), .Q(
        pipeline_regfile_data[242]) );
  DFF_X1 pipeline_regfile_data_reg_8__18_ ( .D(n5008), .CK(clk), .Q(
        pipeline_regfile_data[274]) );
  DFF_X1 pipeline_regfile_data_reg_9__18_ ( .D(n5009), .CK(clk), .Q(
        pipeline_regfile_data[306]) );
  DFF_X1 pipeline_regfile_data_reg_10__18_ ( .D(n5010), .CK(clk), .Q(
        pipeline_regfile_data[338]) );
  DFF_X1 pipeline_regfile_data_reg_11__18_ ( .D(n5011), .CK(clk), .Q(
        pipeline_regfile_data[370]) );
  DFF_X1 pipeline_regfile_data_reg_12__18_ ( .D(n5012), .CK(clk), .Q(
        pipeline_regfile_data[402]) );
  DFF_X1 pipeline_regfile_data_reg_13__18_ ( .D(n5013), .CK(clk), .Q(
        pipeline_regfile_data[434]) );
  DFF_X1 pipeline_regfile_data_reg_14__18_ ( .D(n5014), .CK(clk), .Q(
        pipeline_regfile_data[466]) );
  DFF_X1 pipeline_regfile_data_reg_15__18_ ( .D(n5015), .CK(clk), .Q(
        pipeline_regfile_data[498]) );
  DFF_X1 pipeline_regfile_data_reg_16__18_ ( .D(n5016), .CK(clk), .Q(
        pipeline_regfile_data[530]) );
  DFF_X1 pipeline_regfile_data_reg_17__18_ ( .D(n5017), .CK(clk), .Q(
        pipeline_regfile_data[562]) );
  DFF_X1 pipeline_regfile_data_reg_18__18_ ( .D(n5018), .CK(clk), .Q(
        pipeline_regfile_data[594]) );
  DFF_X1 pipeline_regfile_data_reg_19__18_ ( .D(n5019), .CK(clk), .Q(
        pipeline_regfile_data[626]) );
  DFF_X1 pipeline_regfile_data_reg_20__18_ ( .D(n5020), .CK(clk), .Q(
        pipeline_regfile_data[658]) );
  DFF_X1 pipeline_regfile_data_reg_21__18_ ( .D(n5021), .CK(clk), .Q(
        pipeline_regfile_data[690]) );
  DFF_X1 pipeline_regfile_data_reg_22__18_ ( .D(n5022), .CK(clk), .Q(
        pipeline_regfile_data[722]) );
  DFF_X1 pipeline_regfile_data_reg_23__18_ ( .D(n5023), .CK(clk), .Q(
        pipeline_regfile_data[754]) );
  DFF_X1 pipeline_regfile_data_reg_24__18_ ( .D(n5024), .CK(clk), .Q(
        pipeline_regfile_data[786]) );
  DFF_X1 pipeline_regfile_data_reg_25__18_ ( .D(n5025), .CK(clk), .Q(
        pipeline_regfile_data[818]) );
  DFF_X1 pipeline_regfile_data_reg_26__18_ ( .D(n5026), .CK(clk), .Q(
        pipeline_regfile_data[850]) );
  DFF_X1 pipeline_regfile_data_reg_27__18_ ( .D(n5027), .CK(clk), .Q(
        pipeline_regfile_data[882]) );
  DFF_X1 pipeline_regfile_data_reg_28__18_ ( .D(n5028), .CK(clk), .Q(
        pipeline_regfile_data[914]) );
  DFF_X1 pipeline_regfile_data_reg_29__18_ ( .D(n5029), .CK(clk), .Q(
        pipeline_regfile_data[946]) );
  DFF_X1 pipeline_regfile_data_reg_30__18_ ( .D(n5030), .CK(clk), .Q(
        pipeline_regfile_data[978]) );
  DFF_X1 pipeline_regfile_data_reg_31__18_ ( .D(n5031), .CK(clk), .Q(
        pipeline_regfile_data[1010]) );
  DFF_X1 pipeline_csr_mtime_full_reg_51_ ( .D(pipeline_csr_N2152), .CK(clk), 
        .Q(pipeline_csr_mtime_full[51]), .QN(n6901) );
  DFF_X1 pipeline_csr_mtime_full_reg_19_ ( .D(pipeline_csr_N2120), .CK(clk), 
        .Q(pipeline_csr_mtime_full[19]) );
  DFF_X1 pipeline_csr_time_full_reg_51_ ( .D(pipeline_csr_N2003), .CK(clk), 
        .Q(pipeline_csr_time_full[51]) );
  DFF_X1 pipeline_csr_time_full_reg_19_ ( .D(pipeline_csr_N1971), .CK(clk), 
        .Q(pipeline_csr_time_full[19]), .QN(n6894) );
  DFF_X1 pipeline_csr_cycle_full_reg_51_ ( .D(pipeline_csr_N1939), .CK(clk), 
        .Q(pipeline_csr_cycle_full[51]) );
  DFF_X1 pipeline_csr_cycle_full_reg_19_ ( .D(pipeline_csr_N1907), .CK(clk), 
        .Q(pipeline_csr_cycle_full[19]) );
  DFF_X1 pipeline_regfile_data_reg_1__19_ ( .D(n4970), .CK(clk), .Q(
        pipeline_regfile_data[51]) );
  DFF_X1 pipeline_regfile_data_reg_2__19_ ( .D(n4971), .CK(clk), .Q(
        pipeline_regfile_data[83]) );
  DFF_X1 pipeline_regfile_data_reg_3__19_ ( .D(n4972), .CK(clk), .Q(
        pipeline_regfile_data[115]) );
  DFF_X1 pipeline_regfile_data_reg_4__19_ ( .D(n4973), .CK(clk), .Q(
        pipeline_regfile_data[147]) );
  DFF_X1 pipeline_regfile_data_reg_5__19_ ( .D(n4974), .CK(clk), .Q(
        pipeline_regfile_data[179]) );
  DFF_X1 pipeline_regfile_data_reg_6__19_ ( .D(n4975), .CK(clk), .Q(
        pipeline_regfile_data[211]) );
  DFF_X1 pipeline_regfile_data_reg_7__19_ ( .D(n4976), .CK(clk), .Q(
        pipeline_regfile_data[243]) );
  DFF_X1 pipeline_regfile_data_reg_8__19_ ( .D(n4977), .CK(clk), .Q(
        pipeline_regfile_data[275]) );
  DFF_X1 pipeline_regfile_data_reg_9__19_ ( .D(n4978), .CK(clk), .Q(
        pipeline_regfile_data[307]) );
  DFF_X1 pipeline_regfile_data_reg_10__19_ ( .D(n4979), .CK(clk), .Q(
        pipeline_regfile_data[339]) );
  DFF_X1 pipeline_regfile_data_reg_11__19_ ( .D(n4980), .CK(clk), .Q(
        pipeline_regfile_data[371]) );
  DFF_X1 pipeline_regfile_data_reg_12__19_ ( .D(n4981), .CK(clk), .Q(
        pipeline_regfile_data[403]) );
  DFF_X1 pipeline_regfile_data_reg_13__19_ ( .D(n4982), .CK(clk), .Q(
        pipeline_regfile_data[435]) );
  DFF_X1 pipeline_regfile_data_reg_14__19_ ( .D(n4983), .CK(clk), .Q(
        pipeline_regfile_data[467]) );
  DFF_X1 pipeline_regfile_data_reg_15__19_ ( .D(n4984), .CK(clk), .Q(
        pipeline_regfile_data[499]) );
  DFF_X1 pipeline_regfile_data_reg_16__19_ ( .D(n4985), .CK(clk), .Q(
        pipeline_regfile_data[531]) );
  DFF_X1 pipeline_regfile_data_reg_17__19_ ( .D(n4986), .CK(clk), .Q(
        pipeline_regfile_data[563]) );
  DFF_X1 pipeline_regfile_data_reg_18__19_ ( .D(n4987), .CK(clk), .Q(
        pipeline_regfile_data[595]) );
  DFF_X1 pipeline_regfile_data_reg_19__19_ ( .D(n4988), .CK(clk), .Q(
        pipeline_regfile_data[627]) );
  DFF_X1 pipeline_regfile_data_reg_20__19_ ( .D(n4989), .CK(clk), .Q(
        pipeline_regfile_data[659]) );
  DFF_X1 pipeline_regfile_data_reg_21__19_ ( .D(n4990), .CK(clk), .Q(
        pipeline_regfile_data[691]) );
  DFF_X1 pipeline_regfile_data_reg_22__19_ ( .D(n4991), .CK(clk), .Q(
        pipeline_regfile_data[723]) );
  DFF_X1 pipeline_regfile_data_reg_23__19_ ( .D(n4992), .CK(clk), .Q(
        pipeline_regfile_data[755]) );
  DFF_X1 pipeline_regfile_data_reg_24__19_ ( .D(n4993), .CK(clk), .Q(
        pipeline_regfile_data[787]) );
  DFF_X1 pipeline_regfile_data_reg_25__19_ ( .D(n4994), .CK(clk), .Q(
        pipeline_regfile_data[819]) );
  DFF_X1 pipeline_regfile_data_reg_26__19_ ( .D(n4995), .CK(clk), .Q(
        pipeline_regfile_data[851]) );
  DFF_X1 pipeline_regfile_data_reg_27__19_ ( .D(n4996), .CK(clk), .Q(
        pipeline_regfile_data[883]) );
  DFF_X1 pipeline_regfile_data_reg_28__19_ ( .D(n4997), .CK(clk), .Q(
        pipeline_regfile_data[915]) );
  DFF_X1 pipeline_regfile_data_reg_29__19_ ( .D(n4998), .CK(clk), .Q(
        pipeline_regfile_data[947]) );
  DFF_X1 pipeline_regfile_data_reg_30__19_ ( .D(n4999), .CK(clk), .Q(
        pipeline_regfile_data[979]) );
  DFF_X1 pipeline_regfile_data_reg_31__19_ ( .D(n5000), .CK(clk), .Q(
        pipeline_regfile_data[1011]) );
  DFF_X2 pipeline_md_b_reg_62_ ( .D(n5718), .CK(clk), .Q(pipeline_md_b[62]), 
        .QN(n1085) );
  DFF_X2 pipeline_md_b_reg_61_ ( .D(n5719), .CK(clk), .Q(pipeline_md_b[61]), 
        .QN(n1084) );
  DFF_X2 pipeline_md_b_reg_60_ ( .D(n5720), .CK(clk), .Q(pipeline_md_b[60]), 
        .QN(n1083) );
  DFF_X2 pipeline_md_b_reg_59_ ( .D(n5721), .CK(clk), .Q(pipeline_md_b[59]), 
        .QN(n1082) );
  DFF_X2 pipeline_md_b_reg_58_ ( .D(n5722), .CK(clk), .Q(pipeline_md_b[58]), 
        .QN(n1081) );
  DFF_X2 pipeline_md_b_reg_57_ ( .D(n5723), .CK(clk), .Q(pipeline_md_b[57]), 
        .QN(n1080) );
  DFF_X2 pipeline_md_b_reg_56_ ( .D(n5724), .CK(clk), .Q(pipeline_md_b[56]), 
        .QN(n1079) );
  DFF_X1 pipeline_csr_mtime_full_reg_52_ ( .D(pipeline_csr_N2153), .CK(clk), 
        .Q(pipeline_csr_mtime_full[52]) );
  DFF_X2 pipeline_csr_instret_full_reg_52_ ( .D(n5994), .CK(clk), .Q(n10889), 
        .QN(n1435) );
  DFF_X1 pipeline_csr_mtime_full_reg_20_ ( .D(pipeline_csr_N2121), .CK(clk), 
        .Q(pipeline_csr_mtime_full[20]), .QN(n6822) );
  DFF_X2 pipeline_csr_time_full_reg_52_ ( .D(pipeline_csr_N2004), .CK(clk), 
        .Q(pipeline_csr_time_full[52]), .QN(n1159) );
  DFF_X1 pipeline_csr_time_full_reg_20_ ( .D(pipeline_csr_N1972), .CK(clk), 
        .Q(pipeline_csr_time_full[20]) );
  DFF_X1 pipeline_csr_cycle_full_reg_52_ ( .D(pipeline_csr_N1940), .CK(clk), 
        .Q(pipeline_csr_cycle_full[52]), .QN(n6880) );
  DFF_X1 pipeline_csr_cycle_full_reg_20_ ( .D(pipeline_csr_N1908), .CK(clk), 
        .Q(pipeline_csr_cycle_full[20]) );
  DFF_X1 pipeline_regfile_data_reg_1__20_ ( .D(n4939), .CK(clk), .Q(
        pipeline_regfile_data[52]) );
  DFF_X1 pipeline_regfile_data_reg_2__20_ ( .D(n4940), .CK(clk), .Q(
        pipeline_regfile_data[84]) );
  DFF_X1 pipeline_regfile_data_reg_3__20_ ( .D(n4941), .CK(clk), .Q(
        pipeline_regfile_data[116]) );
  DFF_X1 pipeline_regfile_data_reg_4__20_ ( .D(n4942), .CK(clk), .Q(
        pipeline_regfile_data[148]) );
  DFF_X1 pipeline_regfile_data_reg_5__20_ ( .D(n4943), .CK(clk), .Q(
        pipeline_regfile_data[180]) );
  DFF_X1 pipeline_regfile_data_reg_6__20_ ( .D(n4944), .CK(clk), .Q(
        pipeline_regfile_data[212]) );
  DFF_X1 pipeline_regfile_data_reg_7__20_ ( .D(n4945), .CK(clk), .Q(
        pipeline_regfile_data[244]) );
  DFF_X1 pipeline_regfile_data_reg_8__20_ ( .D(n4946), .CK(clk), .Q(
        pipeline_regfile_data[276]) );
  DFF_X1 pipeline_regfile_data_reg_9__20_ ( .D(n4947), .CK(clk), .Q(
        pipeline_regfile_data[308]) );
  DFF_X1 pipeline_regfile_data_reg_10__20_ ( .D(n4948), .CK(clk), .Q(
        pipeline_regfile_data[340]) );
  DFF_X1 pipeline_regfile_data_reg_11__20_ ( .D(n4949), .CK(clk), .Q(
        pipeline_regfile_data[372]) );
  DFF_X1 pipeline_regfile_data_reg_12__20_ ( .D(n4950), .CK(clk), .Q(
        pipeline_regfile_data[404]) );
  DFF_X1 pipeline_regfile_data_reg_13__20_ ( .D(n4951), .CK(clk), .Q(
        pipeline_regfile_data[436]) );
  DFF_X1 pipeline_regfile_data_reg_14__20_ ( .D(n4952), .CK(clk), .Q(
        pipeline_regfile_data[468]) );
  DFF_X1 pipeline_regfile_data_reg_15__20_ ( .D(n4953), .CK(clk), .Q(
        pipeline_regfile_data[500]) );
  DFF_X1 pipeline_regfile_data_reg_16__20_ ( .D(n4954), .CK(clk), .Q(
        pipeline_regfile_data[532]) );
  DFF_X1 pipeline_regfile_data_reg_17__20_ ( .D(n4955), .CK(clk), .Q(
        pipeline_regfile_data[564]) );
  DFF_X1 pipeline_regfile_data_reg_18__20_ ( .D(n4956), .CK(clk), .Q(
        pipeline_regfile_data[596]) );
  DFF_X1 pipeline_regfile_data_reg_19__20_ ( .D(n4957), .CK(clk), .Q(
        pipeline_regfile_data[628]) );
  DFF_X1 pipeline_regfile_data_reg_20__20_ ( .D(n4958), .CK(clk), .Q(
        pipeline_regfile_data[660]) );
  DFF_X1 pipeline_regfile_data_reg_21__20_ ( .D(n4959), .CK(clk), .Q(
        pipeline_regfile_data[692]) );
  DFF_X1 pipeline_regfile_data_reg_22__20_ ( .D(n4960), .CK(clk), .Q(
        pipeline_regfile_data[724]) );
  DFF_X1 pipeline_regfile_data_reg_23__20_ ( .D(n4961), .CK(clk), .Q(
        pipeline_regfile_data[756]) );
  DFF_X1 pipeline_regfile_data_reg_24__20_ ( .D(n4962), .CK(clk), .Q(
        pipeline_regfile_data[788]) );
  DFF_X1 pipeline_regfile_data_reg_25__20_ ( .D(n4963), .CK(clk), .Q(
        pipeline_regfile_data[820]) );
  DFF_X1 pipeline_regfile_data_reg_26__20_ ( .D(n4964), .CK(clk), .Q(
        pipeline_regfile_data[852]) );
  DFF_X1 pipeline_regfile_data_reg_27__20_ ( .D(n4965), .CK(clk), .Q(
        pipeline_regfile_data[884]) );
  DFF_X1 pipeline_regfile_data_reg_28__20_ ( .D(n4966), .CK(clk), .Q(
        pipeline_regfile_data[916]) );
  DFF_X1 pipeline_regfile_data_reg_29__20_ ( .D(n4967), .CK(clk), .Q(
        pipeline_regfile_data[948]) );
  DFF_X1 pipeline_regfile_data_reg_30__20_ ( .D(n4968), .CK(clk), .Q(
        pipeline_regfile_data[980]) );
  DFF_X1 pipeline_regfile_data_reg_31__20_ ( .D(n4969), .CK(clk), .Q(
        pipeline_regfile_data[1012]) );
  DFF_X1 pipeline_csr_mtime_full_reg_53_ ( .D(pipeline_csr_N2154), .CK(clk), 
        .Q(pipeline_csr_mtime_full[53]), .QN(n6909) );
  DFF_X1 pipeline_csr_mtime_full_reg_21_ ( .D(pipeline_csr_N2122), .CK(clk), 
        .Q(pipeline_csr_mtime_full[21]) );
  DFF_X1 pipeline_csr_time_full_reg_53_ ( .D(pipeline_csr_N2005), .CK(clk), 
        .Q(pipeline_csr_time_full[53]) );
  DFF_X1 pipeline_csr_time_full_reg_21_ ( .D(pipeline_csr_N1973), .CK(clk), 
        .Q(pipeline_csr_time_full[21]), .QN(n6892) );
  DFF_X1 pipeline_csr_cycle_full_reg_53_ ( .D(pipeline_csr_N1941), .CK(clk), 
        .Q(pipeline_csr_cycle_full[53]) );
  DFF_X1 pipeline_csr_cycle_full_reg_21_ ( .D(pipeline_csr_N1909), .CK(clk), 
        .Q(pipeline_csr_cycle_full[21]) );
  DFF_X1 pipeline_regfile_data_reg_1__21_ ( .D(n4908), .CK(clk), .Q(
        pipeline_regfile_data[53]) );
  DFF_X1 pipeline_regfile_data_reg_2__21_ ( .D(n4909), .CK(clk), .Q(
        pipeline_regfile_data[85]) );
  DFF_X1 pipeline_regfile_data_reg_3__21_ ( .D(n4910), .CK(clk), .Q(
        pipeline_regfile_data[117]) );
  DFF_X1 pipeline_regfile_data_reg_4__21_ ( .D(n4911), .CK(clk), .Q(
        pipeline_regfile_data[149]) );
  DFF_X1 pipeline_regfile_data_reg_5__21_ ( .D(n4912), .CK(clk), .Q(
        pipeline_regfile_data[181]) );
  DFF_X1 pipeline_regfile_data_reg_6__21_ ( .D(n4913), .CK(clk), .Q(
        pipeline_regfile_data[213]) );
  DFF_X1 pipeline_regfile_data_reg_7__21_ ( .D(n4914), .CK(clk), .Q(
        pipeline_regfile_data[245]) );
  DFF_X1 pipeline_regfile_data_reg_8__21_ ( .D(n4915), .CK(clk), .Q(
        pipeline_regfile_data[277]) );
  DFF_X1 pipeline_regfile_data_reg_9__21_ ( .D(n4916), .CK(clk), .Q(
        pipeline_regfile_data[309]) );
  DFF_X1 pipeline_regfile_data_reg_10__21_ ( .D(n4917), .CK(clk), .Q(
        pipeline_regfile_data[341]) );
  DFF_X1 pipeline_regfile_data_reg_11__21_ ( .D(n4918), .CK(clk), .Q(
        pipeline_regfile_data[373]) );
  DFF_X1 pipeline_regfile_data_reg_12__21_ ( .D(n4919), .CK(clk), .Q(
        pipeline_regfile_data[405]) );
  DFF_X1 pipeline_regfile_data_reg_13__21_ ( .D(n4920), .CK(clk), .Q(
        pipeline_regfile_data[437]) );
  DFF_X1 pipeline_regfile_data_reg_14__21_ ( .D(n4921), .CK(clk), .Q(
        pipeline_regfile_data[469]) );
  DFF_X1 pipeline_regfile_data_reg_15__21_ ( .D(n4922), .CK(clk), .Q(
        pipeline_regfile_data[501]) );
  DFF_X1 pipeline_regfile_data_reg_16__21_ ( .D(n4923), .CK(clk), .Q(
        pipeline_regfile_data[533]) );
  DFF_X1 pipeline_regfile_data_reg_17__21_ ( .D(n4924), .CK(clk), .Q(
        pipeline_regfile_data[565]) );
  DFF_X1 pipeline_regfile_data_reg_18__21_ ( .D(n4925), .CK(clk), .Q(
        pipeline_regfile_data[597]) );
  DFF_X1 pipeline_regfile_data_reg_19__21_ ( .D(n4926), .CK(clk), .Q(
        pipeline_regfile_data[629]) );
  DFF_X1 pipeline_regfile_data_reg_20__21_ ( .D(n4927), .CK(clk), .Q(
        pipeline_regfile_data[661]) );
  DFF_X1 pipeline_regfile_data_reg_21__21_ ( .D(n4928), .CK(clk), .Q(
        pipeline_regfile_data[693]) );
  DFF_X1 pipeline_regfile_data_reg_22__21_ ( .D(n4929), .CK(clk), .Q(
        pipeline_regfile_data[725]) );
  DFF_X1 pipeline_regfile_data_reg_23__21_ ( .D(n4930), .CK(clk), .Q(
        pipeline_regfile_data[757]) );
  DFF_X1 pipeline_regfile_data_reg_24__21_ ( .D(n4931), .CK(clk), .Q(
        pipeline_regfile_data[789]) );
  DFF_X1 pipeline_regfile_data_reg_25__21_ ( .D(n4932), .CK(clk), .Q(
        pipeline_regfile_data[821]) );
  DFF_X1 pipeline_regfile_data_reg_26__21_ ( .D(n4933), .CK(clk), .Q(
        pipeline_regfile_data[853]) );
  DFF_X1 pipeline_regfile_data_reg_27__21_ ( .D(n4934), .CK(clk), .Q(
        pipeline_regfile_data[885]) );
  DFF_X1 pipeline_regfile_data_reg_28__21_ ( .D(n4935), .CK(clk), .Q(
        pipeline_regfile_data[917]) );
  DFF_X1 pipeline_regfile_data_reg_29__21_ ( .D(n4936), .CK(clk), .Q(
        pipeline_regfile_data[949]) );
  DFF_X1 pipeline_regfile_data_reg_30__21_ ( .D(n4937), .CK(clk), .Q(
        pipeline_regfile_data[981]) );
  DFF_X1 pipeline_regfile_data_reg_31__21_ ( .D(n4938), .CK(clk), .Q(
        pipeline_regfile_data[1013]) );
  DFF_X1 pipeline_csr_mtime_full_reg_22_ ( .D(pipeline_csr_N2123), .CK(clk), 
        .Q(pipeline_csr_mtime_full[22]) );
  DFF_X1 pipeline_csr_time_full_reg_54_ ( .D(pipeline_csr_N2006), .CK(clk), 
        .Q(pipeline_csr_time_full[54]) );
  DFF_X1 pipeline_csr_time_full_reg_22_ ( .D(pipeline_csr_N1974), .CK(clk), 
        .Q(pipeline_csr_time_full[22]), .QN(n6863) );
  DFF_X1 pipeline_csr_cycle_full_reg_54_ ( .D(pipeline_csr_N1942), .CK(clk), 
        .Q(pipeline_csr_cycle_full[54]) );
  DFF_X1 pipeline_csr_cycle_full_reg_22_ ( .D(pipeline_csr_N1910), .CK(clk), 
        .Q(pipeline_csr_cycle_full[22]) );
  DFF_X1 pipeline_regfile_data_reg_1__22_ ( .D(n4877), .CK(clk), .Q(
        pipeline_regfile_data[54]) );
  DFF_X1 pipeline_regfile_data_reg_2__22_ ( .D(n4878), .CK(clk), .Q(
        pipeline_regfile_data[86]) );
  DFF_X1 pipeline_regfile_data_reg_3__22_ ( .D(n4879), .CK(clk), .Q(
        pipeline_regfile_data[118]) );
  DFF_X1 pipeline_regfile_data_reg_4__22_ ( .D(n4880), .CK(clk), .Q(
        pipeline_regfile_data[150]) );
  DFF_X1 pipeline_regfile_data_reg_5__22_ ( .D(n4881), .CK(clk), .Q(
        pipeline_regfile_data[182]) );
  DFF_X1 pipeline_regfile_data_reg_6__22_ ( .D(n4882), .CK(clk), .Q(
        pipeline_regfile_data[214]) );
  DFF_X1 pipeline_regfile_data_reg_7__22_ ( .D(n4883), .CK(clk), .Q(
        pipeline_regfile_data[246]) );
  DFF_X1 pipeline_regfile_data_reg_8__22_ ( .D(n4884), .CK(clk), .Q(
        pipeline_regfile_data[278]) );
  DFF_X1 pipeline_regfile_data_reg_9__22_ ( .D(n4885), .CK(clk), .Q(
        pipeline_regfile_data[310]) );
  DFF_X1 pipeline_regfile_data_reg_10__22_ ( .D(n4886), .CK(clk), .Q(
        pipeline_regfile_data[342]) );
  DFF_X1 pipeline_regfile_data_reg_11__22_ ( .D(n4887), .CK(clk), .Q(
        pipeline_regfile_data[374]) );
  DFF_X1 pipeline_regfile_data_reg_12__22_ ( .D(n4888), .CK(clk), .Q(
        pipeline_regfile_data[406]) );
  DFF_X1 pipeline_regfile_data_reg_13__22_ ( .D(n4889), .CK(clk), .Q(
        pipeline_regfile_data[438]) );
  DFF_X1 pipeline_regfile_data_reg_14__22_ ( .D(n4890), .CK(clk), .Q(
        pipeline_regfile_data[470]) );
  DFF_X1 pipeline_regfile_data_reg_15__22_ ( .D(n4891), .CK(clk), .Q(
        pipeline_regfile_data[502]) );
  DFF_X1 pipeline_regfile_data_reg_16__22_ ( .D(n4892), .CK(clk), .Q(
        pipeline_regfile_data[534]) );
  DFF_X1 pipeline_regfile_data_reg_17__22_ ( .D(n4893), .CK(clk), .Q(
        pipeline_regfile_data[566]) );
  DFF_X1 pipeline_regfile_data_reg_18__22_ ( .D(n4894), .CK(clk), .Q(
        pipeline_regfile_data[598]) );
  DFF_X1 pipeline_regfile_data_reg_19__22_ ( .D(n4895), .CK(clk), .Q(
        pipeline_regfile_data[630]) );
  DFF_X1 pipeline_regfile_data_reg_20__22_ ( .D(n4896), .CK(clk), .Q(
        pipeline_regfile_data[662]) );
  DFF_X1 pipeline_regfile_data_reg_21__22_ ( .D(n4897), .CK(clk), .Q(
        pipeline_regfile_data[694]) );
  DFF_X1 pipeline_regfile_data_reg_22__22_ ( .D(n4898), .CK(clk), .Q(
        pipeline_regfile_data[726]) );
  DFF_X1 pipeline_regfile_data_reg_23__22_ ( .D(n4899), .CK(clk), .Q(
        pipeline_regfile_data[758]) );
  DFF_X1 pipeline_regfile_data_reg_24__22_ ( .D(n4900), .CK(clk), .Q(
        pipeline_regfile_data[790]) );
  DFF_X1 pipeline_regfile_data_reg_25__22_ ( .D(n4901), .CK(clk), .Q(
        pipeline_regfile_data[822]) );
  DFF_X1 pipeline_regfile_data_reg_26__22_ ( .D(n4902), .CK(clk), .Q(
        pipeline_regfile_data[854]) );
  DFF_X1 pipeline_regfile_data_reg_27__22_ ( .D(n4903), .CK(clk), .Q(
        pipeline_regfile_data[886]) );
  DFF_X1 pipeline_regfile_data_reg_28__22_ ( .D(n4904), .CK(clk), .Q(
        pipeline_regfile_data[918]) );
  DFF_X1 pipeline_regfile_data_reg_29__22_ ( .D(n4905), .CK(clk), .Q(
        pipeline_regfile_data[950]) );
  DFF_X1 pipeline_regfile_data_reg_30__22_ ( .D(n4906), .CK(clk), .Q(
        pipeline_regfile_data[982]) );
  DFF_X1 pipeline_regfile_data_reg_31__22_ ( .D(n4907), .CK(clk), .Q(
        pipeline_regfile_data[1014]) );
  DFF_X1 pipeline_regfile_data_reg_1__23_ ( .D(n4846), .CK(clk), .Q(
        pipeline_regfile_data[55]) );
  DFF_X1 pipeline_regfile_data_reg_2__23_ ( .D(n4847), .CK(clk), .Q(
        pipeline_regfile_data[87]) );
  DFF_X1 pipeline_regfile_data_reg_3__23_ ( .D(n4848), .CK(clk), .Q(
        pipeline_regfile_data[119]) );
  DFF_X1 pipeline_regfile_data_reg_4__23_ ( .D(n4849), .CK(clk), .Q(
        pipeline_regfile_data[151]) );
  DFF_X1 pipeline_regfile_data_reg_5__23_ ( .D(n4850), .CK(clk), .Q(
        pipeline_regfile_data[183]) );
  DFF_X1 pipeline_regfile_data_reg_6__23_ ( .D(n4851), .CK(clk), .Q(
        pipeline_regfile_data[215]) );
  DFF_X1 pipeline_regfile_data_reg_7__23_ ( .D(n4852), .CK(clk), .Q(
        pipeline_regfile_data[247]) );
  DFF_X1 pipeline_regfile_data_reg_8__23_ ( .D(n4853), .CK(clk), .Q(
        pipeline_regfile_data[279]) );
  DFF_X1 pipeline_regfile_data_reg_9__23_ ( .D(n4854), .CK(clk), .Q(
        pipeline_regfile_data[311]) );
  DFF_X1 pipeline_regfile_data_reg_10__23_ ( .D(n4855), .CK(clk), .Q(
        pipeline_regfile_data[343]) );
  DFF_X1 pipeline_regfile_data_reg_11__23_ ( .D(n4856), .CK(clk), .Q(
        pipeline_regfile_data[375]) );
  DFF_X1 pipeline_regfile_data_reg_12__23_ ( .D(n4857), .CK(clk), .Q(
        pipeline_regfile_data[407]) );
  DFF_X1 pipeline_regfile_data_reg_13__23_ ( .D(n4858), .CK(clk), .Q(
        pipeline_regfile_data[439]) );
  DFF_X1 pipeline_regfile_data_reg_14__23_ ( .D(n4859), .CK(clk), .Q(
        pipeline_regfile_data[471]) );
  DFF_X1 pipeline_regfile_data_reg_15__23_ ( .D(n4860), .CK(clk), .Q(
        pipeline_regfile_data[503]) );
  DFF_X1 pipeline_regfile_data_reg_16__23_ ( .D(n4861), .CK(clk), .Q(
        pipeline_regfile_data[535]) );
  DFF_X1 pipeline_regfile_data_reg_17__23_ ( .D(n4862), .CK(clk), .Q(
        pipeline_regfile_data[567]) );
  DFF_X1 pipeline_regfile_data_reg_18__23_ ( .D(n4863), .CK(clk), .Q(
        pipeline_regfile_data[599]) );
  DFF_X1 pipeline_regfile_data_reg_19__23_ ( .D(n4864), .CK(clk), .Q(
        pipeline_regfile_data[631]) );
  DFF_X1 pipeline_regfile_data_reg_20__23_ ( .D(n4865), .CK(clk), .Q(
        pipeline_regfile_data[663]) );
  DFF_X1 pipeline_regfile_data_reg_21__23_ ( .D(n4866), .CK(clk), .Q(
        pipeline_regfile_data[695]) );
  DFF_X1 pipeline_regfile_data_reg_22__23_ ( .D(n4867), .CK(clk), .Q(
        pipeline_regfile_data[727]) );
  DFF_X1 pipeline_regfile_data_reg_23__23_ ( .D(n4868), .CK(clk), .Q(
        pipeline_regfile_data[759]) );
  DFF_X1 pipeline_regfile_data_reg_24__23_ ( .D(n4869), .CK(clk), .Q(
        pipeline_regfile_data[791]) );
  DFF_X1 pipeline_regfile_data_reg_25__23_ ( .D(n4870), .CK(clk), .Q(
        pipeline_regfile_data[823]) );
  DFF_X1 pipeline_regfile_data_reg_26__23_ ( .D(n4871), .CK(clk), .Q(
        pipeline_regfile_data[855]) );
  DFF_X1 pipeline_regfile_data_reg_27__23_ ( .D(n4872), .CK(clk), .Q(
        pipeline_regfile_data[887]) );
  DFF_X1 pipeline_regfile_data_reg_28__23_ ( .D(n4873), .CK(clk), .Q(
        pipeline_regfile_data[919]) );
  DFF_X1 pipeline_regfile_data_reg_29__23_ ( .D(n4874), .CK(clk), .Q(
        pipeline_regfile_data[951]) );
  DFF_X1 pipeline_regfile_data_reg_30__23_ ( .D(n4875), .CK(clk), .Q(
        pipeline_regfile_data[983]) );
  DFF_X1 pipeline_regfile_data_reg_31__23_ ( .D(n4876), .CK(clk), .Q(
        pipeline_regfile_data[1015]) );
  DFF_X2 pipeline_md_a_reg_24_ ( .D(n5676), .CK(clk), .Q(pipeline_md_a[24]), 
        .QN(n1111) );
  DFF_X1 pipeline_regfile_data_reg_1__24_ ( .D(n4815), .CK(clk), .Q(
        pipeline_regfile_data[56]) );
  DFF_X1 pipeline_regfile_data_reg_2__24_ ( .D(n4816), .CK(clk), .Q(
        pipeline_regfile_data[88]) );
  DFF_X1 pipeline_regfile_data_reg_3__24_ ( .D(n4817), .CK(clk), .Q(
        pipeline_regfile_data[120]) );
  DFF_X1 pipeline_regfile_data_reg_4__24_ ( .D(n4818), .CK(clk), .Q(
        pipeline_regfile_data[152]) );
  DFF_X1 pipeline_regfile_data_reg_5__24_ ( .D(n4819), .CK(clk), .Q(
        pipeline_regfile_data[184]) );
  DFF_X1 pipeline_regfile_data_reg_6__24_ ( .D(n4820), .CK(clk), .Q(
        pipeline_regfile_data[216]) );
  DFF_X1 pipeline_regfile_data_reg_7__24_ ( .D(n4821), .CK(clk), .Q(
        pipeline_regfile_data[248]) );
  DFF_X1 pipeline_regfile_data_reg_8__24_ ( .D(n4822), .CK(clk), .Q(
        pipeline_regfile_data[280]) );
  DFF_X1 pipeline_regfile_data_reg_9__24_ ( .D(n4823), .CK(clk), .Q(
        pipeline_regfile_data[312]) );
  DFF_X1 pipeline_regfile_data_reg_10__24_ ( .D(n4824), .CK(clk), .Q(
        pipeline_regfile_data[344]) );
  DFF_X1 pipeline_regfile_data_reg_11__24_ ( .D(n4825), .CK(clk), .Q(
        pipeline_regfile_data[376]) );
  DFF_X1 pipeline_regfile_data_reg_12__24_ ( .D(n4826), .CK(clk), .Q(
        pipeline_regfile_data[408]) );
  DFF_X1 pipeline_regfile_data_reg_13__24_ ( .D(n4827), .CK(clk), .Q(
        pipeline_regfile_data[440]) );
  DFF_X1 pipeline_regfile_data_reg_14__24_ ( .D(n4828), .CK(clk), .Q(
        pipeline_regfile_data[472]) );
  DFF_X1 pipeline_regfile_data_reg_15__24_ ( .D(n4829), .CK(clk), .Q(
        pipeline_regfile_data[504]) );
  DFF_X1 pipeline_regfile_data_reg_16__24_ ( .D(n4830), .CK(clk), .Q(
        pipeline_regfile_data[536]) );
  DFF_X1 pipeline_regfile_data_reg_17__24_ ( .D(n4831), .CK(clk), .Q(
        pipeline_regfile_data[568]) );
  DFF_X1 pipeline_regfile_data_reg_18__24_ ( .D(n4832), .CK(clk), .Q(
        pipeline_regfile_data[600]) );
  DFF_X1 pipeline_regfile_data_reg_19__24_ ( .D(n4833), .CK(clk), .Q(
        pipeline_regfile_data[632]) );
  DFF_X1 pipeline_regfile_data_reg_20__24_ ( .D(n4834), .CK(clk), .Q(
        pipeline_regfile_data[664]) );
  DFF_X1 pipeline_regfile_data_reg_21__24_ ( .D(n4835), .CK(clk), .Q(
        pipeline_regfile_data[696]) );
  DFF_X1 pipeline_regfile_data_reg_22__24_ ( .D(n4836), .CK(clk), .Q(
        pipeline_regfile_data[728]) );
  DFF_X1 pipeline_regfile_data_reg_23__24_ ( .D(n4837), .CK(clk), .Q(
        pipeline_regfile_data[760]) );
  DFF_X1 pipeline_regfile_data_reg_24__24_ ( .D(n4838), .CK(clk), .Q(
        pipeline_regfile_data[792]) );
  DFF_X1 pipeline_regfile_data_reg_25__24_ ( .D(n4839), .CK(clk), .Q(
        pipeline_regfile_data[824]) );
  DFF_X1 pipeline_regfile_data_reg_26__24_ ( .D(n4840), .CK(clk), .Q(
        pipeline_regfile_data[856]) );
  DFF_X1 pipeline_regfile_data_reg_27__24_ ( .D(n4841), .CK(clk), .Q(
        pipeline_regfile_data[888]) );
  DFF_X1 pipeline_regfile_data_reg_28__24_ ( .D(n4842), .CK(clk), .Q(
        pipeline_regfile_data[920]) );
  DFF_X1 pipeline_regfile_data_reg_29__24_ ( .D(n4843), .CK(clk), .Q(
        pipeline_regfile_data[952]) );
  DFF_X1 pipeline_regfile_data_reg_30__24_ ( .D(n4844), .CK(clk), .Q(
        pipeline_regfile_data[984]) );
  DFF_X1 pipeline_regfile_data_reg_31__24_ ( .D(n4845), .CK(clk), .Q(
        pipeline_regfile_data[1016]) );
  DFF_X2 pipeline_md_a_reg_25_ ( .D(n5677), .CK(clk), .Q(pipeline_md_a[25]), 
        .QN(n1112) );
  DFF_X1 pipeline_regfile_data_reg_1__25_ ( .D(n4784), .CK(clk), .Q(
        pipeline_regfile_data[57]) );
  DFF_X1 pipeline_regfile_data_reg_2__25_ ( .D(n4785), .CK(clk), .Q(
        pipeline_regfile_data[89]) );
  DFF_X1 pipeline_regfile_data_reg_3__25_ ( .D(n4786), .CK(clk), .Q(
        pipeline_regfile_data[121]) );
  DFF_X1 pipeline_regfile_data_reg_4__25_ ( .D(n4787), .CK(clk), .Q(
        pipeline_regfile_data[153]) );
  DFF_X1 pipeline_regfile_data_reg_5__25_ ( .D(n4788), .CK(clk), .Q(
        pipeline_regfile_data[185]) );
  DFF_X1 pipeline_regfile_data_reg_6__25_ ( .D(n4789), .CK(clk), .Q(
        pipeline_regfile_data[217]) );
  DFF_X1 pipeline_regfile_data_reg_7__25_ ( .D(n4790), .CK(clk), .Q(
        pipeline_regfile_data[249]) );
  DFF_X1 pipeline_regfile_data_reg_8__25_ ( .D(n4791), .CK(clk), .Q(
        pipeline_regfile_data[281]) );
  DFF_X1 pipeline_regfile_data_reg_9__25_ ( .D(n4792), .CK(clk), .Q(
        pipeline_regfile_data[313]) );
  DFF_X1 pipeline_regfile_data_reg_10__25_ ( .D(n4793), .CK(clk), .Q(
        pipeline_regfile_data[345]) );
  DFF_X1 pipeline_regfile_data_reg_11__25_ ( .D(n4794), .CK(clk), .Q(
        pipeline_regfile_data[377]) );
  DFF_X1 pipeline_regfile_data_reg_12__25_ ( .D(n4795), .CK(clk), .Q(
        pipeline_regfile_data[409]) );
  DFF_X1 pipeline_regfile_data_reg_13__25_ ( .D(n4796), .CK(clk), .Q(
        pipeline_regfile_data[441]) );
  DFF_X1 pipeline_regfile_data_reg_14__25_ ( .D(n4797), .CK(clk), .Q(
        pipeline_regfile_data[473]) );
  DFF_X1 pipeline_regfile_data_reg_15__25_ ( .D(n4798), .CK(clk), .Q(
        pipeline_regfile_data[505]) );
  DFF_X1 pipeline_regfile_data_reg_16__25_ ( .D(n4799), .CK(clk), .Q(
        pipeline_regfile_data[537]) );
  DFF_X1 pipeline_regfile_data_reg_17__25_ ( .D(n4800), .CK(clk), .Q(
        pipeline_regfile_data[569]) );
  DFF_X1 pipeline_regfile_data_reg_18__25_ ( .D(n4801), .CK(clk), .Q(
        pipeline_regfile_data[601]) );
  DFF_X1 pipeline_regfile_data_reg_19__25_ ( .D(n4802), .CK(clk), .Q(
        pipeline_regfile_data[633]) );
  DFF_X1 pipeline_regfile_data_reg_20__25_ ( .D(n4803), .CK(clk), .Q(
        pipeline_regfile_data[665]) );
  DFF_X1 pipeline_regfile_data_reg_21__25_ ( .D(n4804), .CK(clk), .Q(
        pipeline_regfile_data[697]) );
  DFF_X1 pipeline_regfile_data_reg_22__25_ ( .D(n4805), .CK(clk), .Q(
        pipeline_regfile_data[729]) );
  DFF_X1 pipeline_regfile_data_reg_23__25_ ( .D(n4806), .CK(clk), .Q(
        pipeline_regfile_data[761]) );
  DFF_X1 pipeline_regfile_data_reg_24__25_ ( .D(n4807), .CK(clk), .Q(
        pipeline_regfile_data[793]) );
  DFF_X1 pipeline_regfile_data_reg_25__25_ ( .D(n4808), .CK(clk), .Q(
        pipeline_regfile_data[825]) );
  DFF_X1 pipeline_regfile_data_reg_26__25_ ( .D(n4809), .CK(clk), .Q(
        pipeline_regfile_data[857]) );
  DFF_X1 pipeline_regfile_data_reg_27__25_ ( .D(n4810), .CK(clk), .Q(
        pipeline_regfile_data[889]) );
  DFF_X1 pipeline_regfile_data_reg_28__25_ ( .D(n4811), .CK(clk), .Q(
        pipeline_regfile_data[921]) );
  DFF_X1 pipeline_regfile_data_reg_29__25_ ( .D(n4812), .CK(clk), .Q(
        pipeline_regfile_data[953]) );
  DFF_X1 pipeline_regfile_data_reg_30__25_ ( .D(n4813), .CK(clk), .Q(
        pipeline_regfile_data[985]) );
  DFF_X1 pipeline_regfile_data_reg_31__25_ ( .D(n4814), .CK(clk), .Q(
        pipeline_regfile_data[1017]) );
  DFF_X2 pipeline_md_a_reg_26_ ( .D(n5678), .CK(clk), .Q(pipeline_md_a[26]), 
        .QN(n13055) );
  DFF_X1 pipeline_regfile_data_reg_2__26_ ( .D(n4754), .CK(clk), .Q(
        pipeline_regfile_data[90]) );
  DFF_X1 pipeline_regfile_data_reg_3__26_ ( .D(n4755), .CK(clk), .Q(
        pipeline_regfile_data[122]) );
  DFF_X1 pipeline_regfile_data_reg_5__26_ ( .D(n4757), .CK(clk), .Q(
        pipeline_regfile_data[186]) );
  DFF_X1 pipeline_regfile_data_reg_7__26_ ( .D(n4759), .CK(clk), .Q(
        pipeline_regfile_data[250]) );
  DFF_X1 pipeline_regfile_data_reg_8__26_ ( .D(n4760), .CK(clk), .Q(
        pipeline_regfile_data[282]) );
  DFF_X1 pipeline_regfile_data_reg_9__26_ ( .D(n4761), .CK(clk), .Q(
        pipeline_regfile_data[314]) );
  DFF_X1 pipeline_regfile_data_reg_10__26_ ( .D(n4762), .CK(clk), .Q(
        pipeline_regfile_data[346]) );
  DFF_X1 pipeline_regfile_data_reg_11__26_ ( .D(n4763), .CK(clk), .Q(
        pipeline_regfile_data[378]) );
  DFF_X1 pipeline_regfile_data_reg_12__26_ ( .D(n4764), .CK(clk), .Q(
        pipeline_regfile_data[410]) );
  DFF_X1 pipeline_regfile_data_reg_13__26_ ( .D(n4765), .CK(clk), .Q(
        pipeline_regfile_data[442]) );
  DFF_X1 pipeline_regfile_data_reg_14__26_ ( .D(n4766), .CK(clk), .Q(
        pipeline_regfile_data[474]) );
  DFF_X1 pipeline_regfile_data_reg_15__26_ ( .D(n4767), .CK(clk), .Q(
        pipeline_regfile_data[506]) );
  DFF_X1 pipeline_regfile_data_reg_16__26_ ( .D(n4768), .CK(clk), .Q(
        pipeline_regfile_data[538]) );
  DFF_X1 pipeline_regfile_data_reg_17__26_ ( .D(n4769), .CK(clk), .Q(
        pipeline_regfile_data[570]) );
  DFF_X1 pipeline_regfile_data_reg_18__26_ ( .D(n4770), .CK(clk), .Q(
        pipeline_regfile_data[602]) );
  DFF_X1 pipeline_regfile_data_reg_19__26_ ( .D(n4771), .CK(clk), .Q(
        pipeline_regfile_data[634]) );
  DFF_X1 pipeline_regfile_data_reg_20__26_ ( .D(n4772), .CK(clk), .Q(
        pipeline_regfile_data[666]) );
  DFF_X1 pipeline_regfile_data_reg_21__26_ ( .D(n4773), .CK(clk), .Q(
        pipeline_regfile_data[698]) );
  DFF_X1 pipeline_regfile_data_reg_22__26_ ( .D(n4774), .CK(clk), .Q(
        pipeline_regfile_data[730]) );
  DFF_X1 pipeline_regfile_data_reg_23__26_ ( .D(n4775), .CK(clk), .Q(
        pipeline_regfile_data[762]) );
  DFF_X1 pipeline_regfile_data_reg_24__26_ ( .D(n4776), .CK(clk), .Q(
        pipeline_regfile_data[794]) );
  DFF_X1 pipeline_regfile_data_reg_25__26_ ( .D(n4777), .CK(clk), .Q(
        pipeline_regfile_data[826]) );
  DFF_X1 pipeline_regfile_data_reg_26__26_ ( .D(n4778), .CK(clk), .Q(
        pipeline_regfile_data[858]) );
  DFF_X1 pipeline_regfile_data_reg_27__26_ ( .D(n4779), .CK(clk), .Q(
        pipeline_regfile_data[890]) );
  DFF_X1 pipeline_regfile_data_reg_28__26_ ( .D(n4780), .CK(clk), .Q(
        pipeline_regfile_data[922]) );
  DFF_X1 pipeline_regfile_data_reg_29__26_ ( .D(n4781), .CK(clk), .Q(
        pipeline_regfile_data[954]) );
  DFF_X1 pipeline_regfile_data_reg_30__26_ ( .D(n4782), .CK(clk), .Q(
        pipeline_regfile_data[986]) );
  DFF_X1 pipeline_regfile_data_reg_31__26_ ( .D(n4783), .CK(clk), .Q(
        pipeline_regfile_data[1018]) );
  DFF_X2 pipeline_md_a_reg_27_ ( .D(n5679), .CK(clk), .Q(pipeline_md_a[27]), 
        .QN(n13054) );
  DFF_X1 pipeline_regfile_data_reg_1__27_ ( .D(n4722), .CK(clk), .Q(
        pipeline_regfile_data[59]) );
  DFF_X1 pipeline_regfile_data_reg_2__27_ ( .D(n4723), .CK(clk), .Q(
        pipeline_regfile_data[91]) );
  DFF_X1 pipeline_regfile_data_reg_3__27_ ( .D(n4724), .CK(clk), .Q(
        pipeline_regfile_data[123]) );
  DFF_X1 pipeline_regfile_data_reg_4__27_ ( .D(n4725), .CK(clk), .Q(
        pipeline_regfile_data[155]) );
  DFF_X1 pipeline_regfile_data_reg_5__27_ ( .D(n4726), .CK(clk), .Q(
        pipeline_regfile_data[187]) );
  DFF_X1 pipeline_regfile_data_reg_6__27_ ( .D(n4727), .CK(clk), .Q(
        pipeline_regfile_data[219]) );
  DFF_X1 pipeline_regfile_data_reg_7__27_ ( .D(n4728), .CK(clk), .Q(
        pipeline_regfile_data[251]) );
  DFF_X1 pipeline_regfile_data_reg_8__27_ ( .D(n4729), .CK(clk), .Q(
        pipeline_regfile_data[283]) );
  DFF_X1 pipeline_regfile_data_reg_9__27_ ( .D(n4730), .CK(clk), .Q(
        pipeline_regfile_data[315]) );
  DFF_X1 pipeline_regfile_data_reg_10__27_ ( .D(n4731), .CK(clk), .Q(
        pipeline_regfile_data[347]) );
  DFF_X1 pipeline_regfile_data_reg_11__27_ ( .D(n4732), .CK(clk), .Q(
        pipeline_regfile_data[379]) );
  DFF_X1 pipeline_regfile_data_reg_12__27_ ( .D(n4733), .CK(clk), .Q(
        pipeline_regfile_data[411]) );
  DFF_X1 pipeline_regfile_data_reg_13__27_ ( .D(n4734), .CK(clk), .Q(
        pipeline_regfile_data[443]) );
  DFF_X1 pipeline_regfile_data_reg_14__27_ ( .D(n4735), .CK(clk), .Q(
        pipeline_regfile_data[475]) );
  DFF_X1 pipeline_regfile_data_reg_15__27_ ( .D(n4736), .CK(clk), .Q(
        pipeline_regfile_data[507]) );
  DFF_X1 pipeline_regfile_data_reg_16__27_ ( .D(n4737), .CK(clk), .Q(
        pipeline_regfile_data[539]) );
  DFF_X1 pipeline_regfile_data_reg_17__27_ ( .D(n4738), .CK(clk), .Q(
        pipeline_regfile_data[571]) );
  DFF_X1 pipeline_regfile_data_reg_18__27_ ( .D(n4739), .CK(clk), .Q(
        pipeline_regfile_data[603]) );
  DFF_X1 pipeline_regfile_data_reg_19__27_ ( .D(n4740), .CK(clk), .Q(
        pipeline_regfile_data[635]) );
  DFF_X1 pipeline_regfile_data_reg_20__27_ ( .D(n4741), .CK(clk), .Q(
        pipeline_regfile_data[667]) );
  DFF_X1 pipeline_regfile_data_reg_21__27_ ( .D(n4742), .CK(clk), .Q(
        pipeline_regfile_data[699]) );
  DFF_X1 pipeline_regfile_data_reg_22__27_ ( .D(n4743), .CK(clk), .Q(
        pipeline_regfile_data[731]) );
  DFF_X1 pipeline_regfile_data_reg_23__27_ ( .D(n4744), .CK(clk), .Q(
        pipeline_regfile_data[763]) );
  DFF_X1 pipeline_regfile_data_reg_24__27_ ( .D(n4745), .CK(clk), .Q(
        pipeline_regfile_data[795]) );
  DFF_X1 pipeline_regfile_data_reg_25__27_ ( .D(n4746), .CK(clk), .Q(
        pipeline_regfile_data[827]) );
  DFF_X1 pipeline_regfile_data_reg_26__27_ ( .D(n4747), .CK(clk), .Q(
        pipeline_regfile_data[859]) );
  DFF_X1 pipeline_regfile_data_reg_27__27_ ( .D(n4748), .CK(clk), .Q(
        pipeline_regfile_data[891]) );
  DFF_X1 pipeline_regfile_data_reg_28__27_ ( .D(n4749), .CK(clk), .Q(
        pipeline_regfile_data[923]) );
  DFF_X1 pipeline_regfile_data_reg_29__27_ ( .D(n4750), .CK(clk), .Q(
        pipeline_regfile_data[955]) );
  DFF_X1 pipeline_regfile_data_reg_30__27_ ( .D(n4751), .CK(clk), .Q(
        pipeline_regfile_data[987]) );
  DFF_X1 pipeline_regfile_data_reg_31__27_ ( .D(n4752), .CK(clk), .Q(
        pipeline_regfile_data[1019]) );
  DFF_X1 pipeline_csr_mtime_full_reg_60_ ( .D(pipeline_csr_N2161), .CK(clk), 
        .Q(pipeline_csr_mtime_full[60]) );
  DFF_X1 pipeline_csr_mtime_full_reg_61_ ( .D(pipeline_csr_N2162), .CK(clk), 
        .Q(pipeline_csr_mtime_full[61]), .QN(n6867) );
  DFF_X1 pipeline_csr_mtime_full_reg_62_ ( .D(pipeline_csr_N2163), .CK(clk), 
        .Q(pipeline_csr_mtime_full[62]), .QN(n6911) );
  DFF_X1 pipeline_csr_mtime_full_reg_63_ ( .D(pipeline_csr_N2164), .CK(clk), 
        .Q(pipeline_csr_mtime_full[63]), .QN(n6846) );
  DFF_X1 pipeline_csr_time_full_reg_29_ ( .D(pipeline_csr_N1981), .CK(clk), 
        .Q(pipeline_csr_time_full[29]), .QN(n6887) );
  DFF_X1 pipeline_csr_cycle_full_reg_61_ ( .D(pipeline_csr_N1949), .CK(clk), 
        .Q(pipeline_csr_cycle_full[61]) );
  DFF_X1 pipeline_csr_cycle_full_reg_29_ ( .D(pipeline_csr_N1917), .CK(clk), 
        .Q(pipeline_csr_cycle_full[29]) );
  DFF_X1 pipeline_csr_time_full_reg_62_ ( .D(pipeline_csr_N2014), .CK(clk), 
        .Q(pipeline_csr_time_full[62]) );
  DFF_X1 pipeline_csr_time_full_reg_63_ ( .D(pipeline_csr_N2015), .CK(clk), 
        .Q(pipeline_csr_time_full[63]), .QN(n6915) );
  DFF_X1 pipeline_csr_cycle_full_reg_30_ ( .D(pipeline_csr_N1918), .CK(clk), 
        .Q(pipeline_csr_cycle_full[30]) );
  DFF_X1 pipeline_csr_cycle_full_reg_63_ ( .D(pipeline_csr_N1951), .CK(clk), 
        .Q(pipeline_csr_cycle_full[63]), .QN(n6758) );
  DFF_X2 pipeline_csr_mtvec_reg_7_ ( .D(n6201), .CK(clk), .Q(n10673), .QN(
        n1198) );
  DFF_X2 pipeline_md_a_reg_28_ ( .D(n5680), .CK(clk), .Q(pipeline_md_a[28]), 
        .QN(n1115) );
  DFF_X1 pipeline_regfile_data_reg_8__28_ ( .D(n4698), .CK(clk), .Q(
        pipeline_regfile_data[284]) );
  DFF_X1 pipeline_regfile_data_reg_9__28_ ( .D(n4699), .CK(clk), .Q(
        pipeline_regfile_data[316]) );
  DFF_X1 pipeline_regfile_data_reg_10__28_ ( .D(n4700), .CK(clk), .Q(
        pipeline_regfile_data[348]) );
  DFF_X1 pipeline_regfile_data_reg_11__28_ ( .D(n4701), .CK(clk), .Q(
        pipeline_regfile_data[380]) );
  DFF_X1 pipeline_regfile_data_reg_12__28_ ( .D(n4702), .CK(clk), .Q(
        pipeline_regfile_data[412]) );
  DFF_X1 pipeline_regfile_data_reg_13__28_ ( .D(n4703), .CK(clk), .Q(
        pipeline_regfile_data[444]) );
  DFF_X1 pipeline_regfile_data_reg_14__28_ ( .D(n4704), .CK(clk), .Q(
        pipeline_regfile_data[476]) );
  DFF_X1 pipeline_regfile_data_reg_15__28_ ( .D(n4705), .CK(clk), .Q(
        pipeline_regfile_data[508]) );
  DFF_X1 pipeline_regfile_data_reg_16__28_ ( .D(n4706), .CK(clk), .Q(
        pipeline_regfile_data[540]) );
  DFF_X1 pipeline_regfile_data_reg_17__28_ ( .D(n4707), .CK(clk), .Q(
        pipeline_regfile_data[572]) );
  DFF_X1 pipeline_regfile_data_reg_18__28_ ( .D(n4708), .CK(clk), .Q(
        pipeline_regfile_data[604]) );
  DFF_X1 pipeline_regfile_data_reg_19__28_ ( .D(n4709), .CK(clk), .Q(
        pipeline_regfile_data[636]) );
  DFF_X1 pipeline_regfile_data_reg_20__28_ ( .D(n4710), .CK(clk), .Q(
        pipeline_regfile_data[668]) );
  DFF_X1 pipeline_regfile_data_reg_21__28_ ( .D(n4711), .CK(clk), .Q(
        pipeline_regfile_data[700]) );
  DFF_X1 pipeline_regfile_data_reg_22__28_ ( .D(n4712), .CK(clk), .Q(
        pipeline_regfile_data[732]) );
  DFF_X1 pipeline_regfile_data_reg_23__28_ ( .D(n4713), .CK(clk), .Q(
        pipeline_regfile_data[764]) );
  DFF_X1 pipeline_regfile_data_reg_24__28_ ( .D(n4714), .CK(clk), .Q(
        pipeline_regfile_data[796]) );
  DFF_X1 pipeline_regfile_data_reg_25__28_ ( .D(n4715), .CK(clk), .Q(
        pipeline_regfile_data[828]) );
  DFF_X1 pipeline_regfile_data_reg_26__28_ ( .D(n4716), .CK(clk), .Q(
        pipeline_regfile_data[860]) );
  DFF_X1 pipeline_regfile_data_reg_27__28_ ( .D(n4717), .CK(clk), .Q(
        pipeline_regfile_data[892]) );
  DFF_X1 pipeline_regfile_data_reg_28__28_ ( .D(n4718), .CK(clk), .Q(
        pipeline_regfile_data[924]) );
  DFF_X1 pipeline_regfile_data_reg_29__28_ ( .D(n4719), .CK(clk), .Q(
        pipeline_regfile_data[956]) );
  DFF_X1 pipeline_regfile_data_reg_30__28_ ( .D(n4720), .CK(clk), .Q(
        pipeline_regfile_data[988]) );
  DFF_X1 pipeline_regfile_data_reg_31__28_ ( .D(n4721), .CK(clk), .Q(
        pipeline_regfile_data[1020]) );
  DFF_X2 pipeline_md_result_reg_61_ ( .D(n5592), .CK(clk), .Q(
        pipeline_md_result[61]), .QN(n956) );
  DFF_X2 pipeline_md_a_reg_29_ ( .D(n5682), .CK(clk), .Q(pipeline_md_a[29]), 
        .QN(n1116) );
  DFF_X1 pipeline_regfile_data_reg_8__29_ ( .D(n4667), .CK(clk), .Q(
        pipeline_regfile_data[285]) );
  DFF_X1 pipeline_regfile_data_reg_9__29_ ( .D(n4668), .CK(clk), .Q(
        pipeline_regfile_data[317]) );
  DFF_X1 pipeline_regfile_data_reg_10__29_ ( .D(n4669), .CK(clk), .Q(
        pipeline_regfile_data[349]) );
  DFF_X1 pipeline_regfile_data_reg_11__29_ ( .D(n4670), .CK(clk), .Q(
        pipeline_regfile_data[381]) );
  DFF_X1 pipeline_regfile_data_reg_12__29_ ( .D(n4671), .CK(clk), .Q(
        pipeline_regfile_data[413]) );
  DFF_X1 pipeline_regfile_data_reg_13__29_ ( .D(n4672), .CK(clk), .Q(
        pipeline_regfile_data[445]) );
  DFF_X1 pipeline_regfile_data_reg_14__29_ ( .D(n4673), .CK(clk), .Q(
        pipeline_regfile_data[477]) );
  DFF_X1 pipeline_regfile_data_reg_15__29_ ( .D(n4674), .CK(clk), .Q(
        pipeline_regfile_data[509]) );
  DFF_X1 pipeline_regfile_data_reg_16__29_ ( .D(n4675), .CK(clk), .Q(
        pipeline_regfile_data[541]) );
  DFF_X1 pipeline_regfile_data_reg_17__29_ ( .D(n4676), .CK(clk), .Q(
        pipeline_regfile_data[573]) );
  DFF_X1 pipeline_regfile_data_reg_18__29_ ( .D(n4677), .CK(clk), .Q(
        pipeline_regfile_data[605]) );
  DFF_X1 pipeline_regfile_data_reg_19__29_ ( .D(n4678), .CK(clk), .Q(
        pipeline_regfile_data[637]) );
  DFF_X1 pipeline_regfile_data_reg_20__29_ ( .D(n4679), .CK(clk), .Q(
        pipeline_regfile_data[669]) );
  DFF_X1 pipeline_regfile_data_reg_21__29_ ( .D(n4680), .CK(clk), .Q(
        pipeline_regfile_data[701]) );
  DFF_X1 pipeline_regfile_data_reg_22__29_ ( .D(n4681), .CK(clk), .Q(
        pipeline_regfile_data[733]) );
  DFF_X1 pipeline_regfile_data_reg_23__29_ ( .D(n4682), .CK(clk), .Q(
        pipeline_regfile_data[765]) );
  DFF_X1 pipeline_regfile_data_reg_24__29_ ( .D(n4683), .CK(clk), .Q(
        pipeline_regfile_data[797]) );
  DFF_X1 pipeline_regfile_data_reg_25__29_ ( .D(n4684), .CK(clk), .Q(
        pipeline_regfile_data[829]) );
  DFF_X1 pipeline_regfile_data_reg_26__29_ ( .D(n4685), .CK(clk), .Q(
        pipeline_regfile_data[861]) );
  DFF_X1 pipeline_regfile_data_reg_27__29_ ( .D(n4686), .CK(clk), .Q(
        pipeline_regfile_data[893]) );
  DFF_X1 pipeline_regfile_data_reg_28__29_ ( .D(n4687), .CK(clk), .Q(
        pipeline_regfile_data[925]) );
  DFF_X1 pipeline_regfile_data_reg_29__29_ ( .D(n4688), .CK(clk), .Q(
        pipeline_regfile_data[957]) );
  DFF_X1 pipeline_regfile_data_reg_30__29_ ( .D(n4689), .CK(clk), .Q(
        pipeline_regfile_data[989]) );
  DFF_X1 pipeline_regfile_data_reg_31__29_ ( .D(n4690), .CK(clk), .Q(
        pipeline_regfile_data[1021]) );
  DFF_X1 pipeline_regfile_data_reg_8__30_ ( .D(n4636), .CK(clk), .Q(
        pipeline_regfile_data[286]) );
  DFF_X1 pipeline_regfile_data_reg_9__30_ ( .D(n4637), .CK(clk), .Q(
        pipeline_regfile_data[318]) );
  DFF_X1 pipeline_regfile_data_reg_10__30_ ( .D(n4638), .CK(clk), .Q(
        pipeline_regfile_data[350]) );
  DFF_X1 pipeline_regfile_data_reg_11__30_ ( .D(n4639), .CK(clk), .Q(
        pipeline_regfile_data[382]) );
  DFF_X1 pipeline_regfile_data_reg_12__30_ ( .D(n4640), .CK(clk), .Q(
        pipeline_regfile_data[414]) );
  DFF_X1 pipeline_regfile_data_reg_13__30_ ( .D(n4641), .CK(clk), .Q(
        pipeline_regfile_data[446]) );
  DFF_X1 pipeline_regfile_data_reg_14__30_ ( .D(n4642), .CK(clk), .Q(
        pipeline_regfile_data[478]) );
  DFF_X1 pipeline_regfile_data_reg_15__30_ ( .D(n4643), .CK(clk), .Q(
        pipeline_regfile_data[510]) );
  DFF_X1 pipeline_regfile_data_reg_16__30_ ( .D(n4644), .CK(clk), .Q(
        pipeline_regfile_data[542]) );
  DFF_X1 pipeline_regfile_data_reg_17__30_ ( .D(n4645), .CK(clk), .Q(
        pipeline_regfile_data[574]) );
  DFF_X1 pipeline_regfile_data_reg_18__30_ ( .D(n4646), .CK(clk), .Q(
        pipeline_regfile_data[606]) );
  DFF_X1 pipeline_regfile_data_reg_19__30_ ( .D(n4647), .CK(clk), .Q(
        pipeline_regfile_data[638]) );
  DFF_X1 pipeline_regfile_data_reg_20__30_ ( .D(n4648), .CK(clk), .Q(
        pipeline_regfile_data[670]) );
  DFF_X1 pipeline_regfile_data_reg_21__30_ ( .D(n4649), .CK(clk), .Q(
        pipeline_regfile_data[702]) );
  DFF_X1 pipeline_regfile_data_reg_22__30_ ( .D(n4650), .CK(clk), .Q(
        pipeline_regfile_data[734]) );
  DFF_X1 pipeline_regfile_data_reg_23__30_ ( .D(n4651), .CK(clk), .Q(
        pipeline_regfile_data[766]) );
  DFF_X1 pipeline_regfile_data_reg_24__30_ ( .D(n4652), .CK(clk), .Q(
        pipeline_regfile_data[798]) );
  DFF_X1 pipeline_regfile_data_reg_25__30_ ( .D(n4653), .CK(clk), .Q(
        pipeline_regfile_data[830]) );
  DFF_X1 pipeline_regfile_data_reg_26__30_ ( .D(n4654), .CK(clk), .Q(
        pipeline_regfile_data[862]) );
  DFF_X1 pipeline_regfile_data_reg_27__30_ ( .D(n4655), .CK(clk), .Q(
        pipeline_regfile_data[894]) );
  DFF_X1 pipeline_regfile_data_reg_28__30_ ( .D(n4656), .CK(clk), .Q(
        pipeline_regfile_data[926]) );
  DFF_X1 pipeline_regfile_data_reg_29__30_ ( .D(n4657), .CK(clk), .Q(
        pipeline_regfile_data[958]) );
  DFF_X1 pipeline_regfile_data_reg_30__30_ ( .D(n4658), .CK(clk), .Q(
        pipeline_regfile_data[990]) );
  DFF_X1 pipeline_regfile_data_reg_31__30_ ( .D(n4659), .CK(clk), .Q(
        pipeline_regfile_data[1022]) );
  DFF_X1 pipeline_regfile_data_reg_8__31_ ( .D(n4605), .CK(clk), .Q(
        pipeline_regfile_data[287]) );
  DFF_X1 pipeline_regfile_data_reg_9__31_ ( .D(n4606), .CK(clk), .Q(
        pipeline_regfile_data[319]) );
  DFF_X1 pipeline_regfile_data_reg_10__31_ ( .D(n4607), .CK(clk), .Q(
        pipeline_regfile_data[351]) );
  DFF_X1 pipeline_regfile_data_reg_11__31_ ( .D(n4608), .CK(clk), .Q(
        pipeline_regfile_data[383]) );
  DFF_X1 pipeline_regfile_data_reg_12__31_ ( .D(n4609), .CK(clk), .Q(
        pipeline_regfile_data[415]) );
  DFF_X1 pipeline_regfile_data_reg_13__31_ ( .D(n4610), .CK(clk), .Q(
        pipeline_regfile_data[447]) );
  DFF_X1 pipeline_regfile_data_reg_14__31_ ( .D(n4611), .CK(clk), .Q(
        pipeline_regfile_data[479]) );
  DFF_X1 pipeline_regfile_data_reg_15__31_ ( .D(n4612), .CK(clk), .Q(
        pipeline_regfile_data[511]) );
  DFF_X1 pipeline_regfile_data_reg_16__31_ ( .D(n4613), .CK(clk), .Q(
        pipeline_regfile_data[543]) );
  DFF_X1 pipeline_regfile_data_reg_17__31_ ( .D(n4614), .CK(clk), .Q(
        pipeline_regfile_data[575]) );
  DFF_X1 pipeline_regfile_data_reg_18__31_ ( .D(n4615), .CK(clk), .Q(
        pipeline_regfile_data[607]) );
  DFF_X1 pipeline_regfile_data_reg_19__31_ ( .D(n4616), .CK(clk), .Q(
        pipeline_regfile_data[639]) );
  DFF_X1 pipeline_regfile_data_reg_20__31_ ( .D(n4617), .CK(clk), .Q(
        pipeline_regfile_data[671]) );
  DFF_X1 pipeline_regfile_data_reg_21__31_ ( .D(n4618), .CK(clk), .Q(
        pipeline_regfile_data[703]) );
  DFF_X1 pipeline_regfile_data_reg_22__31_ ( .D(n4619), .CK(clk), .Q(
        pipeline_regfile_data[735]) );
  DFF_X1 pipeline_regfile_data_reg_23__31_ ( .D(n4620), .CK(clk), .Q(
        pipeline_regfile_data[767]) );
  DFF_X1 pipeline_regfile_data_reg_24__31_ ( .D(n4621), .CK(clk), .Q(
        pipeline_regfile_data[799]) );
  DFF_X1 pipeline_regfile_data_reg_25__31_ ( .D(n4622), .CK(clk), .Q(
        pipeline_regfile_data[831]) );
  DFF_X1 pipeline_regfile_data_reg_26__31_ ( .D(n4623), .CK(clk), .Q(
        pipeline_regfile_data[863]) );
  DFF_X1 pipeline_regfile_data_reg_27__31_ ( .D(n4624), .CK(clk), .Q(
        pipeline_regfile_data[895]) );
  DFF_X1 pipeline_regfile_data_reg_28__31_ ( .D(n4625), .CK(clk), .Q(
        pipeline_regfile_data[927]) );
  DFF_X1 pipeline_regfile_data_reg_29__31_ ( .D(n4626), .CK(clk), .Q(
        pipeline_regfile_data[959]) );
  DFF_X1 pipeline_regfile_data_reg_30__31_ ( .D(n4627), .CK(clk), .Q(
        pipeline_regfile_data[991]) );
  DFF_X1 pipeline_regfile_data_reg_31__31_ ( .D(n4628), .CK(clk), .Q(
        pipeline_regfile_data[1023]) );
  DFF_X1 pipeline_regfile_data_reg_1__0_ ( .D(n5559), .CK(clk), .Q(
        pipeline_regfile_data[32]) );
  DFF_X1 pipeline_regfile_data_reg_2__0_ ( .D(n5560), .CK(clk), .Q(
        pipeline_regfile_data[64]) );
  DFF_X1 pipeline_regfile_data_reg_3__0_ ( .D(n5561), .CK(clk), .Q(
        pipeline_regfile_data[96]) );
  DFF_X1 pipeline_regfile_data_reg_4__0_ ( .D(n5562), .CK(clk), .Q(
        pipeline_regfile_data[128]) );
  DFF_X1 pipeline_regfile_data_reg_5__0_ ( .D(n5563), .CK(clk), .Q(
        pipeline_regfile_data[160]) );
  DFF_X1 pipeline_regfile_data_reg_6__0_ ( .D(n5564), .CK(clk), .Q(
        pipeline_regfile_data[192]) );
  DFF_X1 pipeline_regfile_data_reg_7__0_ ( .D(n5565), .CK(clk), .Q(
        pipeline_regfile_data[224]) );
  DFF_X1 pipeline_regfile_data_reg_8__0_ ( .D(n5566), .CK(clk), .Q(
        pipeline_regfile_data[256]) );
  DFF_X1 pipeline_regfile_data_reg_9__0_ ( .D(n5567), .CK(clk), .Q(
        pipeline_regfile_data[288]) );
  DFF_X1 pipeline_regfile_data_reg_10__0_ ( .D(n5568), .CK(clk), .Q(
        pipeline_regfile_data[320]) );
  DFF_X1 pipeline_regfile_data_reg_11__0_ ( .D(n5569), .CK(clk), .Q(
        pipeline_regfile_data[352]) );
  DFF_X1 pipeline_regfile_data_reg_12__0_ ( .D(n5570), .CK(clk), .Q(
        pipeline_regfile_data[384]) );
  DFF_X1 pipeline_regfile_data_reg_13__0_ ( .D(n5571), .CK(clk), .Q(
        pipeline_regfile_data[416]) );
  DFF_X1 pipeline_regfile_data_reg_14__0_ ( .D(n5572), .CK(clk), .Q(
        pipeline_regfile_data[448]) );
  DFF_X1 pipeline_regfile_data_reg_15__0_ ( .D(n5573), .CK(clk), .Q(
        pipeline_regfile_data[480]) );
  DFF_X1 pipeline_regfile_data_reg_16__0_ ( .D(n5574), .CK(clk), .Q(
        pipeline_regfile_data[512]) );
  DFF_X1 pipeline_regfile_data_reg_17__0_ ( .D(n5575), .CK(clk), .Q(
        pipeline_regfile_data[544]) );
  DFF_X1 pipeline_regfile_data_reg_18__0_ ( .D(n5576), .CK(clk), .Q(
        pipeline_regfile_data[576]) );
  DFF_X1 pipeline_regfile_data_reg_19__0_ ( .D(n5577), .CK(clk), .Q(
        pipeline_regfile_data[608]) );
  DFF_X1 pipeline_regfile_data_reg_20__0_ ( .D(n5578), .CK(clk), .Q(
        pipeline_regfile_data[640]) );
  DFF_X1 pipeline_regfile_data_reg_21__0_ ( .D(n5579), .CK(clk), .Q(
        pipeline_regfile_data[672]) );
  DFF_X1 pipeline_regfile_data_reg_22__0_ ( .D(n5580), .CK(clk), .Q(
        pipeline_regfile_data[704]) );
  DFF_X1 pipeline_regfile_data_reg_23__0_ ( .D(n5581), .CK(clk), .Q(
        pipeline_regfile_data[736]) );
  DFF_X1 pipeline_regfile_data_reg_24__0_ ( .D(n5582), .CK(clk), .Q(
        pipeline_regfile_data[768]) );
  DFF_X1 pipeline_regfile_data_reg_25__0_ ( .D(n5583), .CK(clk), .Q(
        pipeline_regfile_data[800]) );
  DFF_X1 pipeline_regfile_data_reg_26__0_ ( .D(n5584), .CK(clk), .Q(
        pipeline_regfile_data[832]) );
  DFF_X1 pipeline_regfile_data_reg_27__0_ ( .D(n5585), .CK(clk), .Q(
        pipeline_regfile_data[864]) );
  DFF_X1 pipeline_regfile_data_reg_28__0_ ( .D(n5586), .CK(clk), .Q(
        pipeline_regfile_data[896]) );
  DFF_X1 pipeline_regfile_data_reg_29__0_ ( .D(n5587), .CK(clk), .Q(
        pipeline_regfile_data[928]) );
  DFF_X1 pipeline_regfile_data_reg_30__0_ ( .D(n5588), .CK(clk), .Q(
        pipeline_regfile_data[960]) );
  DFF_X1 pipeline_regfile_data_reg_31__0_ ( .D(n5589), .CK(clk), .Q(
        pipeline_regfile_data[992]) );
  NOR4_X2 U100 ( .A1(pipeline_md_N21), .A2(pipeline_md_N22), .A3(n1562), .A4(
        pipeline_md_N23), .ZN(n1558) );
  OAI221_X2 U697 ( .B1(n1254), .B2(n6707), .C1(n1286), .C2(n13138), .A(n2008), 
        .ZN(n4566) );
  NAND2_X2 U698 ( .A1(htif_pcr_resp_data[31]), .A2(n2009), .ZN(n2008) );
  OAI221_X2 U699 ( .B1(n10249), .B2(n6707), .C1(n1285), .C2(n13138), .A(n2010), 
        .ZN(n4567) );
  NAND2_X2 U700 ( .A1(htif_pcr_resp_data[30]), .A2(n9532), .ZN(n2010) );
  OAI221_X2 U701 ( .B1(n10365), .B2(n6707), .C1(n1284), .C2(n13138), .A(n2011), 
        .ZN(n4568) );
  NAND2_X2 U702 ( .A1(htif_pcr_resp_data[29]), .A2(n9532), .ZN(n2011) );
  OAI221_X2 U703 ( .B1(n1251), .B2(n6707), .C1(n1283), .C2(n13138), .A(n2012), 
        .ZN(n4569) );
  NAND2_X2 U704 ( .A1(htif_pcr_resp_data[28]), .A2(n2009), .ZN(n2012) );
  OAI221_X2 U705 ( .B1(n10468), .B2(n6707), .C1(n1282), .C2(n13138), .A(n2013), 
        .ZN(n4570) );
  NAND2_X2 U706 ( .A1(htif_pcr_resp_data[27]), .A2(n2009), .ZN(n2013) );
  OAI221_X2 U707 ( .B1(n10544), .B2(n6707), .C1(n1281), .C2(n13138), .A(n2014), 
        .ZN(n4571) );
  NAND2_X2 U708 ( .A1(htif_pcr_resp_data[26]), .A2(n2009), .ZN(n2014) );
  OAI221_X2 U709 ( .B1(n10598), .B2(n6707), .C1(n1280), .C2(n13138), .A(n2015), 
        .ZN(n4572) );
  NAND2_X2 U710 ( .A1(htif_pcr_resp_data[25]), .A2(n2009), .ZN(n2015) );
  OAI221_X2 U711 ( .B1(n10652), .B2(n6707), .C1(n1279), .C2(n13138), .A(n2016), 
        .ZN(n4573) );
  NAND2_X2 U712 ( .A1(htif_pcr_resp_data[24]), .A2(n2009), .ZN(n2016) );
  OAI221_X2 U713 ( .B1(n10706), .B2(n6707), .C1(n1278), .C2(n13138), .A(n2017), 
        .ZN(n4574) );
  NAND2_X2 U714 ( .A1(htif_pcr_resp_data[23]), .A2(n2009), .ZN(n2017) );
  OAI221_X2 U715 ( .B1(n10757), .B2(n6707), .C1(n1277), .C2(n13138), .A(n2018), 
        .ZN(n4575) );
  NAND2_X2 U716 ( .A1(htif_pcr_resp_data[22]), .A2(n2009), .ZN(n2018) );
  OAI221_X2 U717 ( .B1(n10842), .B2(n6707), .C1(n1276), .C2(n13138), .A(n2019), 
        .ZN(n4576) );
  NAND2_X2 U718 ( .A1(htif_pcr_resp_data[21]), .A2(n2009), .ZN(n2019) );
  OAI221_X2 U719 ( .B1(n1243), .B2(n6707), .C1(n1275), .C2(n13138), .A(n2020), 
        .ZN(n4577) );
  NAND2_X2 U720 ( .A1(htif_pcr_resp_data[20]), .A2(n2009), .ZN(n2020) );
  OAI221_X2 U721 ( .B1(n10950), .B2(n6707), .C1(n1274), .C2(n13138), .A(n2021), 
        .ZN(n4578) );
  NAND2_X2 U722 ( .A1(htif_pcr_resp_data[19]), .A2(n2009), .ZN(n2021) );
  OAI221_X2 U723 ( .B1(n10997), .B2(n6707), .C1(n1273), .C2(n13138), .A(n2022), 
        .ZN(n4579) );
  NAND2_X2 U724 ( .A1(htif_pcr_resp_data[18]), .A2(n2009), .ZN(n2022) );
  OAI221_X2 U725 ( .B1(n11057), .B2(n6707), .C1(n1272), .C2(n13138), .A(n2023), 
        .ZN(n4580) );
  NAND2_X2 U726 ( .A1(htif_pcr_resp_data[17]), .A2(n2009), .ZN(n2023) );
  OAI221_X2 U727 ( .B1(n11084), .B2(n6707), .C1(n1271), .C2(n13138), .A(n2024), 
        .ZN(n4581) );
  NAND2_X2 U728 ( .A1(htif_pcr_resp_data[16]), .A2(n2009), .ZN(n2024) );
  OAI221_X2 U729 ( .B1(n1238), .B2(n6707), .C1(n1270), .C2(n13138), .A(n2025), 
        .ZN(n4582) );
  NAND2_X2 U730 ( .A1(htif_pcr_resp_data[15]), .A2(n2009), .ZN(n2025) );
  OAI221_X2 U731 ( .B1(n11142), .B2(n6707), .C1(n1269), .C2(n13138), .A(n2026), 
        .ZN(n4583) );
  NAND2_X2 U732 ( .A1(htif_pcr_resp_data[14]), .A2(n2009), .ZN(n2026) );
  OAI221_X2 U733 ( .B1(n11030), .B2(n6707), .C1(n1268), .C2(n13138), .A(n2027), 
        .ZN(n4584) );
  NAND2_X2 U734 ( .A1(htif_pcr_resp_data[13]), .A2(n2009), .ZN(n2027) );
  OAI221_X2 U735 ( .B1(n10869), .B2(n6707), .C1(n1267), .C2(n13138), .A(n2028), 
        .ZN(n4585) );
  NAND2_X2 U736 ( .A1(htif_pcr_resp_data[12]), .A2(n2009), .ZN(n2028) );
  OAI221_X2 U737 ( .B1(n10923), .B2(n6707), .C1(n1266), .C2(n13138), .A(n2029), 
        .ZN(n4586) );
  NAND2_X2 U738 ( .A1(htif_pcr_resp_data[11]), .A2(n2009), .ZN(n2029) );
  OAI221_X2 U739 ( .B1(n10977), .B2(n6707), .C1(n1265), .C2(n13138), .A(n2030), 
        .ZN(n4587) );
  NAND2_X2 U740 ( .A1(htif_pcr_resp_data[10]), .A2(n2009), .ZN(n2030) );
  OAI221_X2 U741 ( .B1(n10571), .B2(n6707), .C1(n1264), .C2(n13138), .A(n2031), 
        .ZN(n4588) );
  NAND2_X2 U742 ( .A1(htif_pcr_resp_data[9]), .A2(n2009), .ZN(n2031) );
  OAI221_X2 U743 ( .B1(n1231), .B2(n6707), .C1(n1263), .C2(n13138), .A(n2032), 
        .ZN(n4589) );
  NAND2_X2 U744 ( .A1(htif_pcr_resp_data[8]), .A2(n2009), .ZN(n2032) );
  OAI221_X2 U745 ( .B1(n10680), .B2(n6707), .C1(n1262), .C2(n13138), .A(n2033), 
        .ZN(n4590) );
  NAND2_X2 U746 ( .A1(htif_pcr_resp_data[7]), .A2(n2009), .ZN(n2033) );
  OAI221_X2 U747 ( .B1(n1229), .B2(n6707), .C1(n1261), .C2(n13138), .A(n2034), 
        .ZN(n4591) );
  NAND2_X2 U748 ( .A1(htif_pcr_resp_data[6]), .A2(n2009), .ZN(n2034) );
  OAI221_X2 U749 ( .B1(n1228), .B2(n6707), .C1(n1260), .C2(n13138), .A(n2035), 
        .ZN(n4592) );
  NAND2_X2 U750 ( .A1(htif_pcr_resp_data[5]), .A2(n2009), .ZN(n2035) );
  OAI221_X2 U751 ( .B1(n11234), .B2(n6707), .C1(n1259), .C2(n13138), .A(n2036), 
        .ZN(n4593) );
  NAND2_X2 U752 ( .A1(htif_pcr_resp_data[4]), .A2(n2009), .ZN(n2036) );
  OAI221_X2 U753 ( .B1(n1226), .B2(n6707), .C1(n1258), .C2(n13138), .A(n2037), 
        .ZN(n4594) );
  NAND2_X2 U754 ( .A1(htif_pcr_resp_data[3]), .A2(n2009), .ZN(n2037) );
  OAI221_X2 U755 ( .B1(n10401), .B2(n6707), .C1(n1257), .C2(n13138), .A(n2038), 
        .ZN(n4595) );
  NAND2_X2 U756 ( .A1(htif_pcr_resp_data[2]), .A2(n2009), .ZN(n2038) );
  OAI221_X2 U757 ( .B1(n1224), .B2(n6707), .C1(n1256), .C2(n13138), .A(n2039), 
        .ZN(n4596) );
  NAND2_X2 U758 ( .A1(htif_pcr_resp_data[1]), .A2(n2009), .ZN(n2039) );
  OAI221_X2 U759 ( .B1(n1223), .B2(n6707), .C1(n1255), .C2(n13138), .A(n2040), 
        .ZN(n4597) );
  NAND2_X2 U760 ( .A1(htif_pcr_resp_data[0]), .A2(n2009), .ZN(n2040) );
  OAI22_X2 U3852 ( .A1(n11234), .A2(n3683), .B1(n1905), .B2(n6703), .ZN(n6077)
         );
  OAI22_X2 U3853 ( .A1(n1226), .A2(n3683), .B1(n1907), .B2(n6703), .ZN(n6078)
         );
  OAI22_X2 U3854 ( .A1(n10401), .A2(n3683), .B1(n1909), .B2(n6703), .ZN(n6079)
         );
  OAI22_X2 U3856 ( .A1(n1223), .A2(n3683), .B1(n1915), .B2(n6703), .ZN(n6081)
         );
  OAI22_X2 U3861 ( .A1(n1257), .A2(n6689), .B1(n1909), .B2(n6659), .ZN(n6083)
         );
  OAI22_X2 U3862 ( .A1(n1258), .A2(n6689), .B1(n1907), .B2(n6659), .ZN(n6084)
         );
  OAI22_X2 U3863 ( .A1(n1259), .A2(n6689), .B1(n1905), .B2(n6659), .ZN(n6085)
         );
  OAI22_X2 U3890 ( .A1(n1255), .A2(n6689), .B1(n1915), .B2(n6659), .ZN(n6112)
         );
  OAI22_X2 U3918 ( .A1(n1165), .A2(n9530), .B1(n1905), .B2(n6688), .ZN(n6140)
         );
  OAI22_X2 U3919 ( .A1(n1164), .A2(n9530), .B1(n1907), .B2(n6688), .ZN(n6141)
         );
  OAI22_X2 U3920 ( .A1(n1163), .A2(n9530), .B1(n1909), .B2(n6688), .ZN(n6142)
         );
  OAI22_X2 U3922 ( .A1(n1161), .A2(n9530), .B1(n1915), .B2(n6688), .ZN(n6144)
         );
  OAI22_X2 U3953 ( .A1(n1291), .A2(n9529), .B1(n1905), .B2(n6702), .ZN(n6172)
         );
  OAI22_X2 U3954 ( .A1(n1290), .A2(n9529), .B1(n1907), .B2(n6702), .ZN(n6173)
         );
  OAI22_X2 U3955 ( .A1(n1289), .A2(n9529), .B1(n1909), .B2(n6702), .ZN(n6174)
         );
  OAI22_X2 U3957 ( .A1(n1287), .A2(n9529), .B1(n1915), .B2(n6702), .ZN(n6176)
         );
  NAND2_X2 U4010 ( .A1(htif_pcr_req_data[5]), .A2(n13131), .ZN(n3711) );
  NAND2_X2 U4015 ( .A1(htif_pcr_req_data[6]), .A2(n13131), .ZN(n3715) );
  NAND2_X2 U4021 ( .A1(htif_pcr_req_data[8]), .A2(n13131), .ZN(n3718) );
  NAND2_X2 U4026 ( .A1(htif_pcr_req_data[9]), .A2(n13131), .ZN(n3721) );
  NAND2_X2 U4031 ( .A1(htif_pcr_req_data[10]), .A2(n13131), .ZN(n3724) );
  NAND2_X2 U4036 ( .A1(htif_pcr_req_data[11]), .A2(n13131), .ZN(n3727) );
  NAND2_X2 U4041 ( .A1(htif_pcr_req_data[12]), .A2(n13131), .ZN(n3730) );
  NAND2_X2 U4046 ( .A1(htif_pcr_req_data[13]), .A2(n13131), .ZN(n3733) );
  NAND2_X2 U4051 ( .A1(htif_pcr_req_data[14]), .A2(n13131), .ZN(n3736) );
  NAND2_X2 U4056 ( .A1(htif_pcr_req_data[15]), .A2(n13131), .ZN(n3739) );
  NAND2_X2 U4061 ( .A1(htif_pcr_req_data[16]), .A2(n13131), .ZN(n3742) );
  NAND2_X2 U4066 ( .A1(htif_pcr_req_data[17]), .A2(n13131), .ZN(n3745) );
  NAND2_X2 U4071 ( .A1(htif_pcr_req_data[18]), .A2(n13131), .ZN(n3748) );
  NAND2_X2 U4076 ( .A1(htif_pcr_req_data[19]), .A2(n13131), .ZN(n3751) );
  NAND2_X2 U4081 ( .A1(htif_pcr_req_data[20]), .A2(n13131), .ZN(n3754) );
  NAND2_X2 U4086 ( .A1(htif_pcr_req_data[21]), .A2(n13131), .ZN(n3757) );
  NAND2_X2 U4091 ( .A1(htif_pcr_req_data[22]), .A2(n13131), .ZN(n3760) );
  NAND2_X2 U4618 ( .A1(htif_pcr_req_data[7]), .A2(n13131), .ZN(n4130) );
  NOR4_X2 U4637 ( .A1(n4148), .A2(n4149), .A3(n4150), .A4(n4151), .ZN(n4147)
         );
  XOR2_X2 U4638 ( .A(pipeline_csr_mtimecmp[31]), .B(
        pipeline_csr_mtime_full[31]), .Z(n4151) );
  XOR2_X2 U4639 ( .A(pipeline_csr_mtimecmp[30]), .B(
        pipeline_csr_mtime_full[30]), .Z(n4150) );
  XOR2_X2 U4640 ( .A(pipeline_csr_mtimecmp[29]), .B(
        pipeline_csr_mtime_full[29]), .Z(n4149) );
  XOR2_X2 U4641 ( .A(pipeline_csr_mtimecmp[28]), .B(
        pipeline_csr_mtime_full[28]), .Z(n4148) );
  NAND2_X2 U4704 ( .A1(n4201), .A2(n3704), .ZN(n3785) );
  NAND2_X2 U4705 ( .A1(htif_pcr_req_rw), .A2(n9533), .ZN(n3704) );
  NAND2_X2 U4706 ( .A1(n2041), .A2(n4201), .ZN(n4184) );
  NOR3_X2 U4707 ( .A1(n9532), .A2(htif_pcr_req_addr[0]), .A3(n2042), .ZN(n2041) );
  NAND4_X2 U4708 ( .A1(htif_pcr_req_addr[9]), .A2(htif_pcr_req_addr[8]), .A3(
        n4202), .A4(n4203), .ZN(n2042) );
  NOR4_X2 U4709 ( .A1(n4204), .A2(htif_pcr_req_addr[1]), .A3(
        htif_pcr_req_addr[3]), .A4(htif_pcr_req_addr[2]), .ZN(n4203) );
  AND3_X2 U4710 ( .A1(htif_pcr_req_addr[10]), .A2(n13140), .A3(
        htif_pcr_req_addr[7]), .ZN(n4202) );
  NAND3_X2 U4712 ( .A1(htif_pcr_req_ready), .A2(n13130), .A3(n4205), .ZN(n4206) );
  NAND3_X2 U4713 ( .A1(n9532), .A2(n13130), .A3(n4207), .ZN(n4205) );
  NAND2_X2 U4714 ( .A1(htif_pcr_resp_ready), .A2(htif_pcr_resp_valid), .ZN(
        n4207) );
  OAI22_X2 U4757 ( .A1(n13143), .A2(n512), .B1(n504), .B2(n4229), .ZN(
        dmem_hwdata[9]) );
  OAI22_X2 U4758 ( .A1(n13143), .A2(n511), .B1(n503), .B2(n4229), .ZN(
        dmem_hwdata[8]) );
  NAND2_X2 U4767 ( .A1(n13144), .A2(pipeline_dmem_type_WB[0]), .ZN(n4230) );
  OAI22_X2 U4768 ( .A1(n510), .A2(n4231), .B1(n13144), .B2(n526), .ZN(
        dmem_hwdata[23]) );
  OAI22_X2 U4769 ( .A1(n509), .A2(n4231), .B1(n13144), .B2(n525), .ZN(
        dmem_hwdata[22]) );
  OAI22_X2 U4770 ( .A1(n508), .A2(n4231), .B1(n13144), .B2(n524), .ZN(
        dmem_hwdata[21]) );
  OAI22_X2 U4771 ( .A1(n507), .A2(n4231), .B1(n13144), .B2(n523), .ZN(
        dmem_hwdata[20]) );
  OAI22_X2 U4772 ( .A1(n506), .A2(n4231), .B1(n13144), .B2(n522), .ZN(
        dmem_hwdata[19]) );
  OAI22_X2 U4773 ( .A1(n505), .A2(n4231), .B1(n13144), .B2(n521), .ZN(
        dmem_hwdata[18]) );
  OAI22_X2 U4774 ( .A1(n504), .A2(n4231), .B1(n13144), .B2(n520), .ZN(
        dmem_hwdata[17]) );
  OAI22_X2 U4775 ( .A1(n503), .A2(n4231), .B1(n13144), .B2(n519), .ZN(
        dmem_hwdata[16]) );
  OAI22_X2 U4776 ( .A1(n13143), .A2(n518), .B1(n510), .B2(n4229), .ZN(
        dmem_hwdata[15]) );
  OAI22_X2 U4777 ( .A1(n13143), .A2(n517), .B1(n509), .B2(n4229), .ZN(
        dmem_hwdata[14]) );
  OAI22_X2 U4778 ( .A1(n13143), .A2(n516), .B1(n508), .B2(n4229), .ZN(
        dmem_hwdata[13]) );
  OAI22_X2 U4779 ( .A1(n13143), .A2(n515), .B1(n507), .B2(n4229), .ZN(
        dmem_hwdata[12]) );
  OAI22_X2 U4780 ( .A1(n13143), .A2(n514), .B1(n506), .B2(n4229), .ZN(
        dmem_hwdata[11]) );
  OAI22_X2 U4781 ( .A1(n13143), .A2(n513), .B1(n505), .B2(n4229), .ZN(
        dmem_hwdata[10]) );
  NAND2_X2 U4783 ( .A1(n12847), .A2(n12848), .ZN(n4231) );
  OR2_X1 U6023 ( .A1(pipeline_md_N25), .A2(pipeline_md_N24), .ZN(n1562) );
  OR3_X1 U6074 ( .A1(htif_pcr_req_addr[6]), .A2(htif_pcr_req_addr[5]), .A3(
        htif_pcr_req_addr[4]), .ZN(n4204) );
  NOR2_X2 U5 ( .A1(pipeline_md_N21), .A2(pipeline_md_N22), .ZN(n143) );
  NOR2_X2 U6 ( .A1(n13128), .A2(pipeline_md_N22), .ZN(n142) );
  OAI22_X2 U29 ( .A1(n152), .A2(n13126), .B1(pipeline_md_N25), .B2(n151), .ZN(
        pipeline_md_N185) );
  DFF_X2 pipeline_inst_DX_reg_14_ ( .D(n6277), .CK(clk), .Q(
        pipeline_dmem_type_2_), .QN(n603) );
  DFF_X2 pipeline_inst_DX_reg_30_ ( .D(n6293), .CK(clk), .Q(
        pipeline_inst_DX[30]), .QN(n713) );
  DFF_X2 pipeline_inst_DX_reg_17_ ( .D(n6280), .CK(clk), .Q(
        pipeline_regfile_N14), .QN(n638) );
  DFF_X2 pipeline_inst_DX_reg_15_ ( .D(n6278), .CK(clk), .Q(
        pipeline_regfile_N12), .QN(n636) );
  DFF_X2 pipeline_PC_IF_reg_0_ ( .D(n5971), .CK(clk), .QN(n12539) );
  DFF_X2 pipeline_PC_DX_reg_27_ ( .D(n5885), .CK(clk), .Q(pipeline_PC_DX[27]), 
        .QN(n742) );
  DFF_X2 pipeline_PC_DX_reg_26_ ( .D(n5887), .CK(clk), .Q(pipeline_PC_DX[26]), 
        .QN(n741) );
  DFF_X2 pipeline_PC_DX_reg_24_ ( .D(n5891), .CK(clk), .Q(pipeline_PC_DX[24]), 
        .QN(n739) );
  DFF_X2 pipeline_PC_DX_reg_23_ ( .D(n5893), .CK(clk), .Q(pipeline_PC_DX[23]), 
        .QN(n738) );
  DFF_X2 pipeline_PC_DX_reg_22_ ( .D(n5895), .CK(clk), .Q(pipeline_PC_DX[22]), 
        .QN(n737) );
  DFF_X2 pipeline_PC_DX_reg_21_ ( .D(n5897), .CK(clk), .Q(pipeline_PC_DX[21]), 
        .QN(n736) );
  DFF_X2 pipeline_PC_DX_reg_20_ ( .D(n5899), .CK(clk), .Q(pipeline_PC_DX[20]), 
        .QN(n735) );
  DFF_X2 pipeline_PC_DX_reg_17_ ( .D(n5905), .CK(clk), .Q(pipeline_PC_DX[17]), 
        .QN(n732) );
  DFF_X2 pipeline_PC_DX_reg_29_ ( .D(n5881), .CK(clk), .Q(pipeline_PC_DX[29]), 
        .QN(n744) );
  DFF_X2 pipeline_PC_DX_reg_28_ ( .D(n5883), .CK(clk), .Q(pipeline_PC_DX[28]), 
        .QN(n743) );
  DFF_X2 pipeline_PC_DX_reg_25_ ( .D(n5889), .CK(clk), .Q(pipeline_PC_DX[25]), 
        .QN(n740) );
  DFF_X2 pipeline_PC_DX_reg_19_ ( .D(n5901), .CK(clk), .Q(pipeline_PC_DX[19]), 
        .QN(n734) );
  DFF_X2 pipeline_PC_DX_reg_18_ ( .D(n5903), .CK(clk), .Q(pipeline_PC_DX[18]), 
        .QN(n733) );
  DFF_X2 pipeline_PC_DX_reg_3_ ( .D(n5933), .CK(clk), .Q(pipeline_PC_DX[3]), 
        .QN(n718) );
  DFF_X2 pipeline_PC_DX_reg_2_ ( .D(n5935), .CK(clk), .Q(pipeline_PC_DX[2]), 
        .QN(n717) );
  DFF_X2 pipeline_inst_DX_reg_11_ ( .D(n6271), .CK(clk), .Q(
        pipeline_inst_DX[11]), .QN(n598) );
  DFF_X2 pipeline_inst_DX_reg_10_ ( .D(n6269), .CK(clk), .Q(
        pipeline_inst_DX[10]), .QN(n597) );
  DFF_X2 pipeline_alu_out_WB_reg_28_ ( .D(n5816), .CK(clk), .Q(
        pipeline_alu_out_WB[28]), .QN(n499) );
  DFF_X2 pipeline_inst_DX_reg_9_ ( .D(n6267), .CK(clk), .Q(pipeline_inst_DX[9]), .QN(n596) );
  DFF_X2 pipeline_PC_DX_reg_4_ ( .D(n5931), .CK(clk), .Q(pipeline_PC_DX[4]), 
        .QN(n719) );
  DFF_X2 pipeline_inst_DX_reg_21_ ( .D(n6284), .CK(clk), .Q(
        pipeline_regfile_N18), .QN(n700) );
  DFF_X2 pipeline_inst_DX_reg_16_ ( .D(n6279), .CK(clk), .Q(
        pipeline_regfile_N13), .QN(n637) );
  DFF_X2 pipeline_inst_DX_reg_22_ ( .D(n6285), .CK(clk), .Q(
        pipeline_regfile_N19), .QN(n702) );
  DFF_X2 pipeline_inst_DX_reg_13_ ( .D(n6275), .CK(clk), .Q(dmem_hsize[1]), 
        .QN(n602) );
  DFF_X2 pipeline_inst_DX_reg_12_ ( .D(n6273), .CK(clk), .Q(dmem_hsize[0]), 
        .QN(n601) );
  DFF_X2 pipeline_inst_DX_reg_20_ ( .D(n6283), .CK(clk), .Q(
        pipeline_regfile_N17), .QN(n693) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_31_ ( .D(n4566), .CK(clk), .Q(
        htif_pcr_resp_data[31]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_30_ ( .D(n4567), .CK(clk), .Q(
        htif_pcr_resp_data[30]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_29_ ( .D(n4568), .CK(clk), .Q(
        htif_pcr_resp_data[29]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_28_ ( .D(n4569), .CK(clk), .Q(
        htif_pcr_resp_data[28]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_27_ ( .D(n4570), .CK(clk), .Q(
        htif_pcr_resp_data[27]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_26_ ( .D(n4571), .CK(clk), .Q(
        htif_pcr_resp_data[26]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_25_ ( .D(n4572), .CK(clk), .Q(
        htif_pcr_resp_data[25]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_24_ ( .D(n4573), .CK(clk), .Q(
        htif_pcr_resp_data[24]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_23_ ( .D(n4574), .CK(clk), .Q(
        htif_pcr_resp_data[23]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_22_ ( .D(n4575), .CK(clk), .Q(
        htif_pcr_resp_data[22]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_21_ ( .D(n4576), .CK(clk), .Q(
        htif_pcr_resp_data[21]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_19_ ( .D(n4578), .CK(clk), .Q(
        htif_pcr_resp_data[19]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_18_ ( .D(n4579), .CK(clk), .Q(
        htif_pcr_resp_data[18]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_17_ ( .D(n4580), .CK(clk), .Q(
        htif_pcr_resp_data[17]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_16_ ( .D(n4581), .CK(clk), .Q(
        htif_pcr_resp_data[16]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_14_ ( .D(n4583), .CK(clk), .Q(
        htif_pcr_resp_data[14]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_13_ ( .D(n4584), .CK(clk), .Q(
        htif_pcr_resp_data[13]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_12_ ( .D(n4585), .CK(clk), .Q(
        htif_pcr_resp_data[12]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_11_ ( .D(n4586), .CK(clk), .Q(
        htif_pcr_resp_data[11]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_10_ ( .D(n4587), .CK(clk), .Q(
        htif_pcr_resp_data[10]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_9_ ( .D(n4588), .CK(clk), .Q(
        htif_pcr_resp_data[9]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_7_ ( .D(n4590), .CK(clk), .Q(
        htif_pcr_resp_data[7]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_5_ ( .D(n4592), .CK(clk), .Q(
        htif_pcr_resp_data[5]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_4_ ( .D(n4593), .CK(clk), .Q(
        htif_pcr_resp_data[4]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_3_ ( .D(n4594), .CK(clk), .Q(
        htif_pcr_resp_data[3]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_2_ ( .D(n4595), .CK(clk), .Q(
        htif_pcr_resp_data[2]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_0_ ( .D(n4597), .CK(clk), .Q(
        htif_pcr_resp_data[0]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_6_ ( .D(n4591), .CK(clk), .Q(
        htif_pcr_resp_data[6]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_1_ ( .D(n4596), .CK(clk), .Q(
        htif_pcr_resp_data[1]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_20_ ( .D(n4577), .CK(clk), .Q(
        htif_pcr_resp_data[20]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_15_ ( .D(n4582), .CK(clk), .Q(
        htif_pcr_resp_data[15]) );
  DFF_X2 pipeline_csr_htif_resp_data_reg_8_ ( .D(n4589), .CK(clk), .Q(
        htif_pcr_resp_data[8]) );
  DFF_X2 pipeline_md_counter_reg_0_ ( .D(n6249), .CK(clk), .Q(pipeline_md_N21), 
        .QN(n13128) );
  DFF_X2 pipeline_md_counter_reg_4_ ( .D(n6246), .CK(clk), .Q(pipeline_md_N25), 
        .QN(n13126) );
  DFF_X2 pipeline_md_counter_reg_3_ ( .D(n6247), .CK(clk), .Q(pipeline_md_N24), 
        .QN(n13145) );
  DFF_X2 pipeline_md_counter_reg_2_ ( .D(n6248), .CK(clk), .Q(pipeline_md_N23), 
        .QN(n13127) );
  DFF_X2 pipeline_regfile_data_reg_0__31_ ( .D(pipeline_regfile_data[31]), 
        .CK(clk), .Q(pipeline_regfile_data[31]) );
  DFF_X2 pipeline_regfile_data_reg_0__30_ ( .D(pipeline_regfile_data[30]), 
        .CK(clk), .Q(pipeline_regfile_data[30]) );
  DFF_X2 pipeline_regfile_data_reg_0__29_ ( .D(pipeline_regfile_data[29]), 
        .CK(clk), .Q(pipeline_regfile_data[29]) );
  DFF_X2 pipeline_regfile_data_reg_0__28_ ( .D(pipeline_regfile_data[28]), 
        .CK(clk), .Q(pipeline_regfile_data[28]) );
  DFF_X2 pipeline_regfile_data_reg_0__27_ ( .D(pipeline_regfile_data[27]), 
        .CK(clk), .Q(pipeline_regfile_data[27]) );
  DFF_X2 pipeline_regfile_data_reg_0__26_ ( .D(pipeline_regfile_data[26]), 
        .CK(clk), .Q(pipeline_regfile_data[26]) );
  DFF_X2 pipeline_regfile_data_reg_0__25_ ( .D(pipeline_regfile_data[25]), 
        .CK(clk), .Q(pipeline_regfile_data[25]) );
  DFF_X2 pipeline_regfile_data_reg_0__24_ ( .D(pipeline_regfile_data[24]), 
        .CK(clk), .Q(pipeline_regfile_data[24]) );
  DFF_X2 pipeline_regfile_data_reg_0__23_ ( .D(pipeline_regfile_data[23]), 
        .CK(clk), .Q(pipeline_regfile_data[23]) );
  DFF_X2 pipeline_regfile_data_reg_0__22_ ( .D(pipeline_regfile_data[22]), 
        .CK(clk), .Q(pipeline_regfile_data[22]) );
  DFF_X2 pipeline_regfile_data_reg_0__21_ ( .D(pipeline_regfile_data[21]), 
        .CK(clk), .Q(pipeline_regfile_data[21]) );
  DFF_X2 pipeline_regfile_data_reg_0__20_ ( .D(pipeline_regfile_data[20]), 
        .CK(clk), .Q(pipeline_regfile_data[20]) );
  DFF_X2 pipeline_regfile_data_reg_0__19_ ( .D(pipeline_regfile_data[19]), 
        .CK(clk), .Q(pipeline_regfile_data[19]) );
  DFF_X2 pipeline_regfile_data_reg_0__18_ ( .D(pipeline_regfile_data[18]), 
        .CK(clk), .Q(pipeline_regfile_data[18]) );
  DFF_X2 pipeline_regfile_data_reg_0__17_ ( .D(pipeline_regfile_data[17]), 
        .CK(clk), .Q(pipeline_regfile_data[17]) );
  DFF_X2 pipeline_regfile_data_reg_0__16_ ( .D(pipeline_regfile_data[16]), 
        .CK(clk), .Q(pipeline_regfile_data[16]) );
  DFF_X2 pipeline_regfile_data_reg_0__15_ ( .D(pipeline_regfile_data[15]), 
        .CK(clk), .Q(pipeline_regfile_data[15]) );
  DFF_X2 pipeline_regfile_data_reg_0__14_ ( .D(pipeline_regfile_data[14]), 
        .CK(clk), .Q(pipeline_regfile_data[14]) );
  DFF_X2 pipeline_regfile_data_reg_0__13_ ( .D(pipeline_regfile_data[13]), 
        .CK(clk), .Q(pipeline_regfile_data[13]) );
  DFF_X2 pipeline_regfile_data_reg_0__12_ ( .D(pipeline_regfile_data[12]), 
        .CK(clk), .Q(pipeline_regfile_data[12]) );
  DFF_X2 pipeline_regfile_data_reg_0__11_ ( .D(pipeline_regfile_data[11]), 
        .CK(clk), .Q(pipeline_regfile_data[11]) );
  DFF_X2 pipeline_regfile_data_reg_0__10_ ( .D(pipeline_regfile_data[10]), 
        .CK(clk), .Q(pipeline_regfile_data[10]) );
  DFF_X2 pipeline_regfile_data_reg_0__9_ ( .D(pipeline_regfile_data[9]), .CK(
        clk), .Q(pipeline_regfile_data[9]) );
  DFF_X2 pipeline_regfile_data_reg_0__8_ ( .D(pipeline_regfile_data[8]), .CK(
        clk), .Q(pipeline_regfile_data[8]) );
  DFF_X2 pipeline_regfile_data_reg_0__7_ ( .D(pipeline_regfile_data[7]), .CK(
        clk), .Q(pipeline_regfile_data[7]) );
  DFF_X2 pipeline_regfile_data_reg_0__6_ ( .D(pipeline_regfile_data[6]), .CK(
        clk), .Q(pipeline_regfile_data[6]) );
  DFF_X2 pipeline_regfile_data_reg_0__5_ ( .D(pipeline_regfile_data[5]), .CK(
        clk), .Q(pipeline_regfile_data[5]) );
  DFF_X2 pipeline_regfile_data_reg_0__4_ ( .D(pipeline_regfile_data[4]), .CK(
        clk), .Q(pipeline_regfile_data[4]) );
  DFF_X2 pipeline_regfile_data_reg_0__3_ ( .D(pipeline_regfile_data[3]), .CK(
        clk), .Q(pipeline_regfile_data[3]) );
  DFF_X2 pipeline_regfile_data_reg_0__2_ ( .D(pipeline_regfile_data[2]), .CK(
        clk), .Q(pipeline_regfile_data[2]) );
  DFF_X2 pipeline_regfile_data_reg_0__1_ ( .D(pipeline_regfile_data[1]), .CK(
        clk), .Q(pipeline_regfile_data[1]) );
  DFF_X2 pipeline_regfile_data_reg_0__0_ ( .D(pipeline_regfile_data[0]), .CK(
        clk), .Q(pipeline_regfile_data[0]) );
  DFF_X2 pipeline_ctrl_prev_ex_code_WB_reg_2_ ( .D(n5979), .CK(clk), .QN(
        n11191) );
  DFF_X2 pipeline_regfile_data_reg_6__30_ ( .D(n4634), .CK(clk), .Q(
        pipeline_regfile_data[222]) );
  DFF_X2 pipeline_regfile_data_reg_6__29_ ( .D(n4665), .CK(clk), .Q(
        pipeline_regfile_data[221]) );
  DFF_X2 pipeline_regfile_data_reg_4__30_ ( .D(n4632), .CK(clk), .Q(
        pipeline_regfile_data[158]) );
  DFF_X2 pipeline_regfile_data_reg_4__29_ ( .D(n4663), .CK(clk), .Q(
        pipeline_regfile_data[157]) );
  DFF_X2 pipeline_regfile_data_reg_2__30_ ( .D(n4630), .CK(clk), .Q(
        pipeline_regfile_data[94]) );
  DFF_X2 pipeline_regfile_data_reg_2__29_ ( .D(n4661), .CK(clk), .Q(
        pipeline_regfile_data[93]) );
  DFF_X2 pipeline_regfile_data_reg_7__30_ ( .D(n4635), .CK(clk), .Q(
        pipeline_regfile_data[254]) );
  DFF_X2 pipeline_regfile_data_reg_5__30_ ( .D(n4633), .CK(clk), .Q(
        pipeline_regfile_data[190]) );
  DFF_X2 pipeline_regfile_data_reg_3__30_ ( .D(n4631), .CK(clk), .Q(
        pipeline_regfile_data[126]) );
  DFF_X2 pipeline_regfile_data_reg_1__30_ ( .D(n4629), .CK(clk), .Q(
        pipeline_regfile_data[62]) );
  DFF_X2 pipeline_regfile_data_reg_7__31_ ( .D(n4604), .CK(clk), .Q(
        pipeline_regfile_data[255]) );
  DFF_X2 pipeline_regfile_data_reg_7__28_ ( .D(n4697), .CK(clk), .Q(
        pipeline_regfile_data[252]) );
  DFF_X2 pipeline_regfile_data_reg_5__31_ ( .D(n4602), .CK(clk), .Q(
        pipeline_regfile_data[191]) );
  DFF_X2 pipeline_regfile_data_reg_5__28_ ( .D(n4695), .CK(clk), .Q(
        pipeline_regfile_data[188]) );
  DFF_X2 pipeline_regfile_data_reg_3__31_ ( .D(n4600), .CK(clk), .Q(
        pipeline_regfile_data[127]) );
  DFF_X2 pipeline_regfile_data_reg_3__28_ ( .D(n4693), .CK(clk), .Q(
        pipeline_regfile_data[124]) );
  DFF_X2 pipeline_regfile_data_reg_1__31_ ( .D(n4598), .CK(clk), .Q(
        pipeline_regfile_data[63]) );
  DFF_X2 pipeline_regfile_data_reg_1__28_ ( .D(n4691), .CK(clk), .Q(
        pipeline_regfile_data[60]) );
  DFF_X2 pipeline_regfile_data_reg_6__31_ ( .D(n4603), .CK(clk), .Q(
        pipeline_regfile_data[223]) );
  DFF_X2 pipeline_regfile_data_reg_6__28_ ( .D(n4696), .CK(clk), .Q(
        pipeline_regfile_data[220]) );
  DFF_X2 pipeline_regfile_data_reg_4__31_ ( .D(n4601), .CK(clk), .Q(
        pipeline_regfile_data[159]) );
  DFF_X2 pipeline_regfile_data_reg_4__28_ ( .D(n4694), .CK(clk), .Q(
        pipeline_regfile_data[156]) );
  DFF_X2 pipeline_regfile_data_reg_2__31_ ( .D(n4599), .CK(clk), .Q(
        pipeline_regfile_data[95]) );
  DFF_X2 pipeline_regfile_data_reg_2__28_ ( .D(n4692), .CK(clk), .Q(
        pipeline_regfile_data[92]) );
  DFF_X2 pipeline_regfile_data_reg_7__29_ ( .D(n4666), .CK(clk), .Q(
        pipeline_regfile_data[253]) );
  DFF_X2 pipeline_regfile_data_reg_5__29_ ( .D(n4664), .CK(clk), .Q(
        pipeline_regfile_data[189]) );
  DFF_X2 pipeline_regfile_data_reg_3__29_ ( .D(n4662), .CK(clk), .Q(
        pipeline_regfile_data[125]) );
  DFF_X2 pipeline_regfile_data_reg_1__29_ ( .D(n4660), .CK(clk), .Q(
        pipeline_regfile_data[61]) );
  DFF_X2 pipeline_regfile_data_reg_1__26_ ( .D(n4753), .CK(clk), .Q(
        pipeline_regfile_data[58]) );
  DFF_X2 pipeline_regfile_data_reg_6__26_ ( .D(n4758), .CK(clk), .Q(
        pipeline_regfile_data[218]) );
  DFF_X2 pipeline_regfile_data_reg_4__26_ ( .D(n4756), .CK(clk), .Q(
        pipeline_regfile_data[154]) );
  DFF_X2 pipeline_csr_htif_state_reg ( .D(n6368), .CK(clk), .Q(
        htif_pcr_resp_valid), .QN(htif_pcr_req_ready) );
  DFF_X2 pipeline_ctrl_reg_to_wr_WB_reg_3_ ( .D(n6268), .CK(clk), .Q(n12995), 
        .QN(n12996) );
  DFF_X2 pipeline_ctrl_reg_to_wr_WB_reg_4_ ( .D(n6270), .CK(clk), .Q(n12992), 
        .QN(n12993) );
  DFF_X2 pipeline_PC_WB_reg_31_ ( .D(n5876), .CK(clk), .Q(n12597) );
  DFF_X2 pipeline_PC_WB_reg_7_ ( .D(n5924), .CK(clk), .Q(n10819), .QN(n542) );
  DFF_X2 pipeline_PC_WB_reg_6_ ( .D(n5926), .CK(clk), .Q(n10820), .QN(n541) );
  DFF_X2 pipeline_PC_WB_reg_5_ ( .D(n5928), .CK(clk), .Q(n10822), .QN(n540) );
  DFF_X2 pipeline_PC_WB_reg_4_ ( .D(n5930), .CK(clk), .Q(n12808) );
  DFF_X2 pipeline_PC_WB_reg_30_ ( .D(n5878), .CK(clk), .Q(n10794), .QN(n565)
         );
  DFF_X2 pipeline_PC_WB_reg_8_ ( .D(n5922), .CK(clk), .Q(n10818), .QN(n543) );
  DFF_X2 pipeline_PC_WB_reg_12_ ( .D(n5914), .CK(clk), .Q(n10814), .QN(n547)
         );
  DFF_X2 pipeline_ctrl_reg_to_wr_WB_reg_0_ ( .D(n6262), .CK(clk), .Q(n12990), 
        .QN(n12991) );
  DFF_X2 pipeline_PC_WB_reg_17_ ( .D(n5904), .CK(clk), .Q(n10809), .QN(n552)
         );
  DFF_X2 pipeline_PC_WB_reg_27_ ( .D(n5884), .CK(clk), .Q(n10797), .QN(n562)
         );
  DFF_X2 pipeline_PC_WB_reg_24_ ( .D(n5890), .CK(clk), .Q(n10801), .QN(n559)
         );
  DFF_X2 pipeline_PC_WB_reg_22_ ( .D(n5894), .CK(clk), .Q(n10803), .QN(n557)
         );
  DFF_X2 pipeline_PC_WB_reg_21_ ( .D(n5896), .CK(clk), .Q(n10804), .QN(n556)
         );
  DFF_X2 pipeline_PC_WB_reg_20_ ( .D(n5898), .CK(clk), .Q(n10805), .QN(n555)
         );
  DFF_X2 pipeline_PC_WB_reg_19_ ( .D(n5900), .CK(clk), .Q(n10806), .QN(n554)
         );
  DFF_X2 pipeline_PC_WB_reg_16_ ( .D(n5906), .CK(clk), .Q(n10810), .QN(n551)
         );
  DFF_X2 pipeline_PC_WB_reg_13_ ( .D(n5912), .CK(clk), .Q(n10813), .QN(n548)
         );
  DFF_X2 pipeline_PC_WB_reg_2_ ( .D(n5934), .CK(clk), .Q(n12290) );
  DFF_X2 pipeline_PC_WB_reg_29_ ( .D(n5880), .CK(clk), .Q(n10795), .QN(n564)
         );
  DFF_X2 pipeline_PC_WB_reg_28_ ( .D(n5882), .CK(clk), .Q(n10796), .QN(n563)
         );
  DFF_X2 pipeline_PC_WB_reg_26_ ( .D(n5886), .CK(clk), .Q(n10799), .QN(n561)
         );
  DFF_X2 pipeline_PC_WB_reg_25_ ( .D(n5888), .CK(clk), .Q(n10800), .QN(n560)
         );
  DFF_X2 pipeline_PC_WB_reg_23_ ( .D(n5892), .CK(clk), .Q(n10802), .QN(n558)
         );
  DFF_X2 pipeline_PC_WB_reg_18_ ( .D(n5902), .CK(clk), .Q(n10807), .QN(n553)
         );
  DFF_X2 pipeline_PC_WB_reg_15_ ( .D(n5908), .CK(clk), .Q(n10811), .QN(n550)
         );
  DFF_X2 pipeline_PC_WB_reg_14_ ( .D(n5910), .CK(clk), .Q(n10812), .QN(n549)
         );
  DFF_X2 pipeline_PC_WB_reg_11_ ( .D(n5916), .CK(clk), .Q(n10815), .QN(n546)
         );
  DFF_X2 pipeline_PC_WB_reg_10_ ( .D(n5918), .CK(clk), .Q(n10816), .QN(n545)
         );
  DFF_X2 pipeline_PC_WB_reg_9_ ( .D(n5920), .CK(clk), .Q(n10817), .QN(n544) );
  DFF_X2 pipeline_PC_WB_reg_3_ ( .D(n5932), .CK(clk), .Q(n12144) );
  DFF_X2 pipeline_store_data_WB_reg_4_ ( .D(n6328), .CK(clk), .Q(
        dmem_hwdata[4]), .QN(n507) );
  DFF_X2 pipeline_store_data_WB_reg_5_ ( .D(n6327), .CK(clk), .Q(
        dmem_hwdata[5]), .QN(n508) );
  DFF_X2 pipeline_store_data_WB_reg_0_ ( .D(n6332), .CK(clk), .Q(
        dmem_hwdata[0]), .QN(n503) );
  DFF_X2 pipeline_store_data_WB_reg_2_ ( .D(n6330), .CK(clk), .Q(
        dmem_hwdata[2]), .QN(n505) );
  DFF_X2 pipeline_store_data_WB_reg_6_ ( .D(n6326), .CK(clk), .Q(
        dmem_hwdata[6]), .QN(n509) );
  DFF_X2 pipeline_store_data_WB_reg_7_ ( .D(n6325), .CK(clk), .Q(
        dmem_hwdata[7]), .QN(n510) );
  DFF_X2 pipeline_store_data_WB_reg_3_ ( .D(n6329), .CK(clk), .Q(
        dmem_hwdata[3]), .QN(n506) );
  DFF_X2 pipeline_store_data_WB_reg_1_ ( .D(n6331), .CK(clk), .Q(
        dmem_hwdata[1]), .QN(n504) );
  DFF_X2 pipeline_ctrl_dmem_en_WB_reg ( .D(n6254), .CK(clk), .Q(
        pipeline_ctrl_dmem_en_WB), .QN(n789) );
  DFF_X2 pipeline_md_b_reg_30_ ( .D(n5750), .CK(clk), .Q(pipeline_md_b[30]), 
        .QN(n1053) );
  DFF_X2 pipeline_md_b_reg_29_ ( .D(n5751), .CK(clk), .Q(pipeline_md_b[29]), 
        .QN(n1052) );
  DFF_X2 pipeline_md_b_reg_28_ ( .D(n5752), .CK(clk), .Q(pipeline_md_b[28]), 
        .QN(n1051) );
  DFF_X2 pipeline_md_b_reg_27_ ( .D(n5753), .CK(clk), .Q(pipeline_md_b[27]), 
        .QN(n1050) );
  DFF_X2 pipeline_md_b_reg_26_ ( .D(n5754), .CK(clk), .Q(pipeline_md_b[26]), 
        .QN(n1049) );
  DFF_X2 pipeline_md_b_reg_25_ ( .D(n5755), .CK(clk), .Q(pipeline_md_b[25]), 
        .QN(n1048) );
  DFF_X2 pipeline_md_b_reg_24_ ( .D(n5756), .CK(clk), .Q(pipeline_md_b[24]), 
        .QN(n1047) );
  DFF_X2 pipeline_md_b_reg_23_ ( .D(n5757), .CK(clk), .Q(pipeline_md_b[23]), 
        .QN(n1046) );
  DFF_X2 pipeline_md_b_reg_22_ ( .D(n5758), .CK(clk), .Q(pipeline_md_b[22]), 
        .QN(n1045) );
  DFF_X2 pipeline_md_b_reg_21_ ( .D(n5759), .CK(clk), .Q(pipeline_md_b[21]), 
        .QN(n1044) );
  DFF_X2 pipeline_md_b_reg_20_ ( .D(n5760), .CK(clk), .Q(pipeline_md_b[20]), 
        .QN(n1043) );
  DFF_X2 pipeline_md_b_reg_19_ ( .D(n5761), .CK(clk), .Q(pipeline_md_b[19]), 
        .QN(n1042) );
  DFF_X2 pipeline_md_b_reg_18_ ( .D(n5762), .CK(clk), .Q(pipeline_md_b[18]), 
        .QN(n1041) );
  DFF_X2 pipeline_md_b_reg_17_ ( .D(n5763), .CK(clk), .Q(pipeline_md_b[17]), 
        .QN(n1040) );
  DFF_X2 pipeline_md_b_reg_16_ ( .D(n5764), .CK(clk), .Q(pipeline_md_b[16]), 
        .QN(n1039) );
  DFF_X2 pipeline_md_b_reg_15_ ( .D(n5765), .CK(clk), .Q(pipeline_md_b[15]), 
        .QN(n1038) );
  DFF_X2 pipeline_md_b_reg_14_ ( .D(n5766), .CK(clk), .Q(pipeline_md_b[14]), 
        .QN(n1037) );
  DFF_X2 pipeline_md_b_reg_13_ ( .D(n5767), .CK(clk), .Q(pipeline_md_b[13]), 
        .QN(n1036) );
  DFF_X2 pipeline_md_b_reg_12_ ( .D(n5768), .CK(clk), .Q(pipeline_md_b[12]), 
        .QN(n1035) );
  DFF_X2 pipeline_md_b_reg_11_ ( .D(n5769), .CK(clk), .Q(pipeline_md_b[11]), 
        .QN(n1034) );
  DFF_X2 pipeline_md_b_reg_10_ ( .D(n5770), .CK(clk), .Q(pipeline_md_b[10]), 
        .QN(n1033) );
  DFF_X2 pipeline_md_b_reg_9_ ( .D(n5771), .CK(clk), .Q(pipeline_md_b[9]), 
        .QN(n1032) );
  DFF_X2 pipeline_md_b_reg_8_ ( .D(n5772), .CK(clk), .Q(pipeline_md_b[8]), 
        .QN(n1031) );
  DFF_X2 pipeline_md_negate_output_reg ( .D(n6241), .CK(clk), .Q(n10192), .QN(
        n962) );
  DFF_X2 pipeline_md_b_reg_7_ ( .D(n5773), .CK(clk), .Q(pipeline_md_b[7]), 
        .QN(n1030) );
  DFF_X2 pipeline_md_a_reg_55_ ( .D(n5708), .CK(clk), .Q(pipeline_md_a[55]), 
        .QN(n1142) );
  DFF_X2 pipeline_md_a_reg_54_ ( .D(n5707), .CK(clk), .Q(pipeline_md_a[54]), 
        .QN(n1141) );
  DFF_X2 pipeline_md_a_reg_53_ ( .D(n5706), .CK(clk), .Q(pipeline_md_a[53]), 
        .QN(n1140) );
  DFF_X2 pipeline_md_a_reg_52_ ( .D(n5705), .CK(clk), .Q(pipeline_md_a[52]), 
        .QN(n1139) );
  DFF_X2 pipeline_md_a_reg_51_ ( .D(n5704), .CK(clk), .Q(pipeline_md_a[51]), 
        .QN(n1138) );
  DFF_X2 pipeline_md_a_reg_50_ ( .D(n5703), .CK(clk), .Q(pipeline_md_a[50]), 
        .QN(n1137) );
  DFF_X2 pipeline_md_a_reg_49_ ( .D(n5702), .CK(clk), .Q(pipeline_md_a[49]), 
        .QN(n1136) );
  DFF_X2 pipeline_md_a_reg_48_ ( .D(n5701), .CK(clk), .Q(pipeline_md_a[48]), 
        .QN(n1135) );
  DFF_X2 pipeline_md_a_reg_47_ ( .D(n5700), .CK(clk), .Q(pipeline_md_a[47]), 
        .QN(n1134) );
  DFF_X2 pipeline_md_a_reg_46_ ( .D(n5699), .CK(clk), .Q(pipeline_md_a[46]), 
        .QN(n1133) );
  DFF_X2 pipeline_md_a_reg_45_ ( .D(n5698), .CK(clk), .Q(pipeline_md_a[45]), 
        .QN(n1132) );
  DFF_X2 pipeline_md_a_reg_44_ ( .D(n5697), .CK(clk), .Q(pipeline_md_a[44]), 
        .QN(n1131) );
  DFF_X2 pipeline_md_a_reg_43_ ( .D(n5696), .CK(clk), .Q(pipeline_md_a[43]), 
        .QN(n1130) );
  DFF_X2 pipeline_md_a_reg_42_ ( .D(n5695), .CK(clk), .Q(pipeline_md_a[42]), 
        .QN(n1129) );
  DFF_X2 pipeline_md_a_reg_41_ ( .D(n5694), .CK(clk), .Q(pipeline_md_a[41]), 
        .QN(n1128) );
  DFF_X2 pipeline_md_a_reg_40_ ( .D(n5693), .CK(clk), .Q(pipeline_md_a[40]), 
        .QN(n1127) );
  DFF_X2 pipeline_md_a_reg_39_ ( .D(n5692), .CK(clk), .Q(pipeline_md_a[39]), 
        .QN(n1126) );
  DFF_X2 pipeline_md_a_reg_38_ ( .D(n5691), .CK(clk), .Q(pipeline_md_a[38]), 
        .QN(n1125) );
  DFF_X2 pipeline_md_a_reg_37_ ( .D(n5690), .CK(clk), .Q(pipeline_md_a[37]), 
        .QN(n1124) );
  DFF_X2 pipeline_md_a_reg_36_ ( .D(n5689), .CK(clk), .Q(pipeline_md_a[36]), 
        .QN(n1123) );
  DFF_X2 pipeline_md_a_reg_35_ ( .D(n5688), .CK(clk), .Q(pipeline_md_a[35]), 
        .QN(n1122) );
  DFF_X2 pipeline_md_a_reg_34_ ( .D(n5687), .CK(clk), .Q(pipeline_md_a[34]), 
        .QN(n1121) );
  DFF_X2 pipeline_md_a_reg_33_ ( .D(n5686), .CK(clk), .Q(pipeline_md_a[33]), 
        .QN(n1120) );
  DFF_X2 pipeline_md_a_reg_32_ ( .D(n5685), .CK(clk), .Q(pipeline_md_a[32]), 
        .QN(n1119) );
  DFF_X2 pipeline_md_a_reg_56_ ( .D(n5709), .CK(clk), .Q(pipeline_md_a[56]), 
        .QN(n1143) );
  DFF_X2 pipeline_md_result_reg_56_ ( .D(n5597), .CK(clk), .Q(
        pipeline_md_result[56]), .QN(n946) );
  DFF_X2 pipeline_md_result_reg_55_ ( .D(n5598), .CK(clk), .Q(
        pipeline_md_result[55]), .QN(n944) );
  DFF_X2 pipeline_md_result_reg_54_ ( .D(n5599), .CK(clk), .Q(
        pipeline_md_result[54]), .QN(n942) );
  DFF_X2 pipeline_md_result_reg_53_ ( .D(n5600), .CK(clk), .Q(
        pipeline_md_result[53]), .QN(n940) );
  DFF_X2 pipeline_md_result_reg_52_ ( .D(n5601), .CK(clk), .Q(
        pipeline_md_result[52]), .QN(n938) );
  DFF_X2 pipeline_md_result_reg_51_ ( .D(n5602), .CK(clk), .Q(
        pipeline_md_result[51]), .QN(n936) );
  DFF_X2 pipeline_md_result_reg_50_ ( .D(n5603), .CK(clk), .Q(
        pipeline_md_result[50]), .QN(n934) );
  DFF_X2 pipeline_md_result_reg_49_ ( .D(n5604), .CK(clk), .Q(
        pipeline_md_result[49]), .QN(n932) );
  DFF_X2 pipeline_md_result_reg_48_ ( .D(n5605), .CK(clk), .Q(
        pipeline_md_result[48]), .QN(n930) );
  DFF_X2 pipeline_md_result_reg_47_ ( .D(n5606), .CK(clk), .Q(
        pipeline_md_result[47]), .QN(n928) );
  DFF_X2 pipeline_md_result_reg_46_ ( .D(n5607), .CK(clk), .Q(
        pipeline_md_result[46]), .QN(n926) );
  DFF_X2 pipeline_md_result_reg_45_ ( .D(n5608), .CK(clk), .Q(
        pipeline_md_result[45]), .QN(n924) );
  DFF_X2 pipeline_md_result_reg_44_ ( .D(n5609), .CK(clk), .Q(
        pipeline_md_result[44]), .QN(n922) );
  DFF_X2 pipeline_md_result_reg_43_ ( .D(n5610), .CK(clk), .Q(
        pipeline_md_result[43]), .QN(n920) );
  DFF_X2 pipeline_md_result_reg_42_ ( .D(n5611), .CK(clk), .Q(
        pipeline_md_result[42]), .QN(n918) );
  DFF_X2 pipeline_md_result_reg_41_ ( .D(n5612), .CK(clk), .Q(
        pipeline_md_result[41]), .QN(n916) );
  DFF_X2 pipeline_md_result_reg_40_ ( .D(n5613), .CK(clk), .Q(
        pipeline_md_result[40]), .QN(n914) );
  DFF_X2 pipeline_md_result_reg_39_ ( .D(n5614), .CK(clk), .Q(
        pipeline_md_result[39]), .QN(n912) );
  DFF_X2 pipeline_md_result_reg_38_ ( .D(n5615), .CK(clk), .Q(
        pipeline_md_result[38]), .QN(n910) );
  DFF_X2 pipeline_md_result_reg_37_ ( .D(n5616), .CK(clk), .Q(
        pipeline_md_result[37]), .QN(n908) );
  DFF_X2 pipeline_md_result_reg_36_ ( .D(n5617), .CK(clk), .Q(
        pipeline_md_result[36]), .QN(n906) );
  DFF_X2 pipeline_md_result_reg_35_ ( .D(n5618), .CK(clk), .Q(
        pipeline_md_result[35]), .QN(n904) );
  DFF_X2 pipeline_md_result_reg_34_ ( .D(n5619), .CK(clk), .Q(
        pipeline_md_result[34]), .QN(n902) );
  DFF_X2 pipeline_md_result_reg_33_ ( .D(n5620), .CK(clk), .Q(
        pipeline_md_result[33]), .QN(n900) );
  DFF_X2 pipeline_md_result_reg_32_ ( .D(n5621), .CK(clk), .Q(
        pipeline_md_result[32]), .QN(n898) );
  DFF_X2 pipeline_md_a_reg_1_ ( .D(n5681), .CK(clk), .Q(pipeline_md_a[1]), 
        .QN(n1088) );
  DFF_X2 pipeline_md_result_reg_57_ ( .D(n5596), .CK(clk), .Q(
        pipeline_md_result[57]), .QN(n948) );
  DFF_X2 pipeline_md_a_reg_15_ ( .D(n5667), .CK(clk), .Q(pipeline_md_a[15]), 
        .QN(n13039) );
  DFF_X2 pipeline_md_a_reg_22_ ( .D(n5674), .CK(clk), .Q(pipeline_md_a[22]), 
        .QN(n13067) );
  DFF_X2 pipeline_md_a_reg_21_ ( .D(n5673), .CK(clk), .Q(pipeline_md_a[21]), 
        .QN(n1108) );
  DFF_X2 pipeline_md_a_reg_20_ ( .D(n5672), .CK(clk), .Q(pipeline_md_a[20]), 
        .QN(n1107) );
  DFF_X2 pipeline_md_a_reg_19_ ( .D(n5671), .CK(clk), .Q(pipeline_md_a[19]), 
        .QN(n13063) );
  DFF_X2 pipeline_md_a_reg_18_ ( .D(n5670), .CK(clk), .Q(pipeline_md_a[18]), 
        .QN(n13064) );
  DFF_X2 pipeline_md_a_reg_17_ ( .D(n5669), .CK(clk), .Q(pipeline_md_a[17]), 
        .QN(n1104) );
  DFF_X2 pipeline_md_a_reg_13_ ( .D(n5665), .CK(clk), .Q(pipeline_md_a[13]), 
        .QN(n1100) );
  DFF_X2 pipeline_md_a_reg_9_ ( .D(n5661), .CK(clk), .Q(pipeline_md_a[9]), 
        .QN(n1096) );
  DFF_X2 pipeline_md_a_reg_7_ ( .D(n5659), .CK(clk), .Q(pipeline_md_a[7]), 
        .QN(n13048) );
  DFF_X2 pipeline_md_a_reg_57_ ( .D(n5710), .CK(clk), .Q(pipeline_md_a[57]), 
        .QN(n1144) );
  DFF_X2 pipeline_md_a_reg_14_ ( .D(n5666), .CK(clk), .Q(pipeline_md_a[14]), 
        .QN(n13040) );
  DFF_X2 pipeline_md_a_reg_23_ ( .D(n5675), .CK(clk), .Q(pipeline_md_a[23]), 
        .QN(n13066) );
  DFF_X2 pipeline_md_b_reg_54_ ( .D(n5726), .CK(clk), .Q(pipeline_md_b[54]), 
        .QN(n1077) );
  DFF_X2 pipeline_md_b_reg_53_ ( .D(n5727), .CK(clk), .Q(pipeline_md_b[53]), 
        .QN(n1076) );
  DFF_X2 pipeline_md_b_reg_52_ ( .D(n5728), .CK(clk), .Q(pipeline_md_b[52]), 
        .QN(n1075) );
  DFF_X2 pipeline_md_b_reg_51_ ( .D(n5729), .CK(clk), .Q(pipeline_md_b[51]), 
        .QN(n1074) );
  DFF_X2 pipeline_md_b_reg_50_ ( .D(n5730), .CK(clk), .Q(pipeline_md_b[50]), 
        .QN(n1073) );
  DFF_X2 pipeline_md_b_reg_49_ ( .D(n5731), .CK(clk), .Q(pipeline_md_b[49]), 
        .QN(n1072) );
  DFF_X2 pipeline_md_b_reg_48_ ( .D(n5732), .CK(clk), .Q(pipeline_md_b[48]), 
        .QN(n1071) );
  DFF_X2 pipeline_md_b_reg_47_ ( .D(n5733), .CK(clk), .Q(pipeline_md_b[47]), 
        .QN(n1070) );
  DFF_X2 pipeline_md_b_reg_46_ ( .D(n5734), .CK(clk), .Q(pipeline_md_b[46]), 
        .QN(n1069) );
  DFF_X2 pipeline_md_b_reg_45_ ( .D(n5735), .CK(clk), .Q(pipeline_md_b[45]), 
        .QN(n1068) );
  DFF_X2 pipeline_md_b_reg_44_ ( .D(n5736), .CK(clk), .Q(pipeline_md_b[44]), 
        .QN(n1067) );
  DFF_X2 pipeline_md_b_reg_42_ ( .D(n5738), .CK(clk), .Q(pipeline_md_b[42]), 
        .QN(n1065) );
  DFF_X2 pipeline_md_b_reg_41_ ( .D(n5739), .CK(clk), .Q(pipeline_md_b[41]), 
        .QN(n1064) );
  DFF_X2 pipeline_md_b_reg_40_ ( .D(n5740), .CK(clk), .Q(pipeline_md_b[40]), 
        .QN(n1063) );
  DFF_X2 pipeline_md_b_reg_37_ ( .D(n5743), .CK(clk), .Q(pipeline_md_b[37]), 
        .QN(n1060) );
  DFF_X2 pipeline_md_b_reg_31_ ( .D(n5749), .CK(clk), .Q(pipeline_md_b[31]), 
        .QN(n1054) );
  DFF_X2 pipeline_csr_mtvec_reg_30_ ( .D(n6178), .CK(clk), .Q(n10238), .QN(
        n1221) );
  DFF_X2 pipeline_csr_mtvec_reg_29_ ( .D(n6179), .CK(clk), .Q(n10358), .QN(
        n1220) );
  DFF_X2 pipeline_csr_mtvec_reg_27_ ( .D(n6181), .CK(clk), .Q(n10461), .QN(
        n1218) );
  DFF_X2 pipeline_csr_mtvec_reg_26_ ( .D(n6182), .CK(clk), .Q(n10537), .QN(
        n1217) );
  DFF_X2 pipeline_csr_mtvec_reg_25_ ( .D(n6183), .CK(clk), .Q(n10591), .QN(
        n1216) );
  DFF_X2 pipeline_csr_mtvec_reg_24_ ( .D(n6184), .CK(clk), .Q(n10645), .QN(
        n1215) );
  DFF_X2 pipeline_csr_mtvec_reg_23_ ( .D(n6185), .CK(clk), .Q(n10699), .QN(
        n1214) );
  DFF_X2 pipeline_csr_mtvec_reg_22_ ( .D(n6186), .CK(clk), .Q(n10750), .QN(
        n1213) );
  DFF_X2 pipeline_csr_mtvec_reg_21_ ( .D(n6187), .CK(clk), .Q(n10835), .QN(
        n1212) );
  DFF_X2 pipeline_csr_mtvec_reg_20_ ( .D(n6188), .CK(clk), .Q(n10895), .QN(
        n1211) );
  DFF_X2 pipeline_csr_mtvec_reg_19_ ( .D(n6189), .CK(clk), .Q(n10943), .QN(
        n1210) );
  DFF_X2 pipeline_csr_mtvec_reg_18_ ( .D(n6190), .CK(clk), .Q(n11003), .QN(
        n1209) );
  DFF_X2 pipeline_csr_mtvec_reg_17_ ( .D(n6191), .CK(clk), .Q(n11050), .QN(
        n1208) );
  DFF_X2 pipeline_csr_mtvec_reg_16_ ( .D(n6192), .CK(clk), .Q(n11077), .QN(
        n1207) );
  DFF_X2 pipeline_csr_mtvec_reg_15_ ( .D(n6193), .CK(clk), .Q(n11113), .QN(
        n1206) );
  DFF_X2 pipeline_csr_mtvec_reg_14_ ( .D(n6194), .CK(clk), .Q(n11133), .QN(
        n1205) );
  DFF_X2 pipeline_csr_mtvec_reg_13_ ( .D(n6195), .CK(clk), .Q(n11023), .QN(
        n1204) );
  DFF_X2 pipeline_csr_mtvec_reg_12_ ( .D(n6196), .CK(clk), .Q(n10862), .QN(
        n1203) );
  DFF_X2 pipeline_csr_mtvec_reg_11_ ( .D(n6197), .CK(clk), .Q(n10916), .QN(
        n1202) );
  DFF_X2 pipeline_csr_mtvec_reg_10_ ( .D(n6198), .CK(clk), .Q(n10970), .QN(
        n1201) );
  DFF_X2 pipeline_csr_mtvec_reg_9_ ( .D(n6199), .CK(clk), .Q(n10564), .QN(
        n1200) );
  DFF_X2 pipeline_csr_mtvec_reg_28_ ( .D(n6180), .CK(clk), .Q(n10426), .QN(
        n1219) );
  DFF_X2 pipeline_md_a_reg_16_ ( .D(n5668), .CK(clk), .Q(pipeline_md_a[16]), 
        .QN(n1103) );
  DFF_X2 pipeline_md_a_reg_12_ ( .D(n5664), .CK(clk), .Q(pipeline_md_a[12]), 
        .QN(n1099) );
  DFF_X2 pipeline_md_a_reg_11_ ( .D(n5663), .CK(clk), .Q(pipeline_md_a[11]), 
        .QN(n13036) );
  DFF_X2 pipeline_md_a_reg_10_ ( .D(n5662), .CK(clk), .Q(pipeline_md_a[10]), 
        .QN(n13037) );
  DFF_X2 pipeline_md_a_reg_8_ ( .D(n5660), .CK(clk), .Q(pipeline_md_a[8]), 
        .QN(n1095) );
  DFF_X2 pipeline_md_a_reg_6_ ( .D(n5658), .CK(clk), .Q(pipeline_md_a[6]), 
        .QN(n13049) );
  DFF_X2 pipeline_md_a_reg_5_ ( .D(n5657), .CK(clk), .Q(pipeline_md_a[5]), 
        .QN(n1092) );
  DFF_X2 pipeline_md_a_reg_3_ ( .D(n5655), .CK(clk), .Q(pipeline_md_a[3]), 
        .QN(n13045) );
  DFF_X2 pipeline_md_a_reg_2_ ( .D(n5654), .CK(clk), .Q(pipeline_md_a[2]), 
        .QN(n13046) );
  DFF_X2 pipeline_md_a_reg_0_ ( .D(n5716), .CK(clk), .Q(pipeline_md_a[0]), 
        .QN(n1087) );
  DFF_X2 pipeline_md_a_reg_4_ ( .D(n5656), .CK(clk), .Q(pipeline_md_a[4]), 
        .QN(n1091) );
  DFF_X2 pipeline_md_b_reg_55_ ( .D(n5725), .CK(clk), .Q(pipeline_md_b[55]), 
        .QN(n1078) );
  DFF_X2 pipeline_md_b_reg_43_ ( .D(n5737), .CK(clk), .Q(pipeline_md_b[43]), 
        .QN(n1066) );
  DFF_X2 pipeline_md_b_reg_39_ ( .D(n5741), .CK(clk), .Q(pipeline_md_b[39]), 
        .QN(n1062) );
  DFF_X2 pipeline_md_b_reg_38_ ( .D(n5742), .CK(clk), .Q(pipeline_md_b[38]), 
        .QN(n1061) );
  DFF_X2 pipeline_md_b_reg_36_ ( .D(n5744), .CK(clk), .Q(pipeline_md_b[36]), 
        .QN(n1059) );
  DFF_X2 pipeline_md_b_reg_35_ ( .D(n5745), .CK(clk), .Q(pipeline_md_b[35]), 
        .QN(n1058) );
  DFF_X2 pipeline_md_b_reg_34_ ( .D(n5746), .CK(clk), .Q(pipeline_md_b[34]), 
        .QN(n1057) );
  DFF_X2 pipeline_md_b_reg_33_ ( .D(n5747), .CK(clk), .Q(pipeline_md_b[33]), 
        .QN(n1056) );
  DFF_X2 pipeline_md_b_reg_32_ ( .D(n5748), .CK(clk), .Q(pipeline_md_b[32]), 
        .QN(n1055) );
  DFF_X2 pipeline_csr_time_full_reg_47_ ( .D(pipeline_csr_N1999), .CK(clk), 
        .Q(pipeline_csr_time_full[47]), .QN(n1158) );
  DFF_X2 pipeline_PC_DX_reg_16_ ( .D(n5907), .CK(clk), .Q(pipeline_PC_DX[16]), 
        .QN(n731) );
  DFF_X2 pipeline_PC_DX_reg_15_ ( .D(n5909), .CK(clk), .Q(pipeline_PC_DX[15]), 
        .QN(n730) );
  DFF_X2 pipeline_PC_DX_reg_14_ ( .D(n5911), .CK(clk), .Q(pipeline_PC_DX[14]), 
        .QN(n729) );
  DFF_X2 pipeline_PC_DX_reg_13_ ( .D(n5913), .CK(clk), .Q(pipeline_PC_DX[13]), 
        .QN(n728) );
  DFF_X2 pipeline_PC_DX_reg_12_ ( .D(n5915), .CK(clk), .Q(pipeline_PC_DX[12]), 
        .QN(n727) );
  DFF_X2 pipeline_PC_DX_reg_11_ ( .D(n5917), .CK(clk), .Q(pipeline_PC_DX[11]), 
        .QN(n726) );
  DFF_X2 pipeline_PC_DX_reg_10_ ( .D(n5919), .CK(clk), .Q(pipeline_PC_DX[10]), 
        .QN(n725) );
  DFF_X2 pipeline_PC_DX_reg_9_ ( .D(n5921), .CK(clk), .Q(pipeline_PC_DX[9]), 
        .QN(n724) );
  DFF_X2 pipeline_alu_out_WB_reg_29_ ( .D(n5815), .CK(clk), .Q(
        pipeline_alu_out_WB[29]), .QN(n500) );
  DFF_X2 pipeline_md_a_reg_63_ ( .D(n5717), .CK(clk), .Q(n10233), .QN(n1150)
         );
  DFF_X2 pipeline_md_result_reg_62_ ( .D(n5591), .CK(clk), .Q(
        pipeline_md_result[62]), .QN(n958) );
  DFF_X2 pipeline_PC_IF_reg_4_ ( .D(n5967), .CK(clk), .QN(n12525) );
  DFF_X2 pipeline_PC_IF_reg_2_ ( .D(n5969), .CK(clk), .QN(n12534) );
  DFF_X2 pipeline_alu_out_WB_reg_31_ ( .D(n5813), .CK(clk), .Q(
        pipeline_alu_out_WB[31]), .QN(n502) );
  DFF_X2 pipeline_PC_IF_reg_16_ ( .D(n5955), .CK(clk), .QN(n12476) );
  DFF_X2 pipeline_md_a_reg_62_ ( .D(n5715), .CK(clk), .Q(pipeline_md_a[62]), 
        .QN(n1149) );
  DFF_X2 pipeline_PC_IF_reg_3_ ( .D(n5968), .CK(clk), .QN(n12529) );
  DFF_X2 pipeline_md_result_reg_63_ ( .D(n5590), .CK(clk), .Q(n10234), .QN(
        n960) );
  DFF_X2 pipeline_PC_IF_reg_12_ ( .D(n5959), .CK(clk), .QN(n12492) );
  DFF_X2 pipeline_PC_IF_reg_13_ ( .D(n5958), .CK(clk), .QN(n12488) );
  DFF_X2 pipeline_PC_IF_reg_17_ ( .D(n5954), .CK(clk), .QN(n12473) );
  DFF_X2 pipeline_PC_IF_reg_5_ ( .D(n5966), .CK(clk), .QN(n12520) );
  DFF_X2 pipeline_PC_IF_reg_15_ ( .D(n5956), .CK(clk), .QN(n12480) );
  DFF_X2 pipeline_PC_IF_reg_8_ ( .D(n5963), .CK(clk), .Q(pipeline_PC_IF_8_), 
        .QN(n12508) );
  DFF_X2 pipeline_alu_out_WB_reg_30_ ( .D(n5814), .CK(clk), .Q(
        pipeline_alu_out_WB[30]), .QN(n501) );
  DFF_X2 pipeline_PC_IF_reg_14_ ( .D(n5957), .CK(clk), .QN(n12484) );
  DFF_X2 pipeline_PC_IF_reg_11_ ( .D(n5960), .CK(clk), .QN(n12496) );
  DFF_X2 pipeline_PC_IF_reg_6_ ( .D(n5965), .CK(clk), .QN(n12516) );
  DFF_X2 pipeline_PC_IF_reg_7_ ( .D(n5964), .CK(clk), .QN(n12512) );
  DFF_X2 pipeline_md_state_reg_1_ ( .D(pipeline_md_N162), .CK(clk), .Q(
        pipeline_md_state[1]), .QN(n9642) );
  DFF_X2 pipeline_ctrl_reg_to_wr_WB_reg_2_ ( .D(n6266), .CK(clk), .Q(
        pipeline_reg_to_wr_WB[2]), .QN(n12988) );
  DFF_X2 pipeline_dmem_type_WB_reg_2_ ( .D(n6276), .CK(clk), .Q(
        pipeline_dmem_type_WB[2]), .QN(n12848) );
  DFF_X2 pipeline_dmem_type_WB_reg_1_ ( .D(n6274), .CK(clk), .Q(
        pipeline_dmem_type_WB[1]), .QN(n12847) );
  DFF_X2 pipeline_dmem_type_WB_reg_0_ ( .D(n6272), .CK(clk), .Q(
        pipeline_dmem_type_WB[0]), .QN(n12846) );
  DFF_X2 pipeline_ctrl_reg_to_wr_WB_reg_1_ ( .D(n6264), .CK(clk), .Q(
        pipeline_reg_to_wr_WB[1]), .QN(n12989) );
  DFF_X2 pipeline_ctrl_wb_src_sel_WB_reg_1_ ( .D(n6333), .CK(clk), .Q(n10144), 
        .QN(n9535) );
  DFF_X2 pipeline_ctrl_wb_src_sel_WB_reg_0_ ( .D(n6255), .CK(clk), .Q(
        pipeline_wb_src_sel_WB_0_), .QN(n784) );
  DFF_X2 pipeline_store_data_WB_reg_31_ ( .D(n13136), .CK(clk), .Q(
        pipeline_store_data_WB_31_), .QN(n534) );
  DFF_X2 pipeline_ctrl_prev_ex_code_WB_reg_3_ ( .D(n5978), .CK(clk), .Q(
        pipeline_ctrl_prev_ex_code_WB[3]) );
  DFF_X2 pipeline_regfile_data_reg_25__3_ ( .D(n5490), .CK(clk), .Q(
        pipeline_regfile_data[803]), .QN(n6935) );
  DFF_X2 pipeline_regfile_data_reg_17__3_ ( .D(n5482), .CK(clk), .Q(
        pipeline_regfile_data[547]), .QN(n6934) );
  DFF_X2 pipeline_regfile_data_reg_19__4_ ( .D(n5453), .CK(clk), .Q(
        pipeline_regfile_data[612]), .QN(n6937) );
  DFF_X2 pipeline_ctrl_prev_ex_code_WB_reg_0_ ( .D(n5977), .CK(clk), .Q(
        pipeline_ctrl_prev_ex_code_WB[0]), .QN(n780) );
  DFF_X2 pipeline_ctrl_had_ex_WB_reg ( .D(n6299), .CK(clk), .Q(
        pipeline_ctrl_had_ex_WB) );
  DFF_X2 pipeline_ctrl_prev_ex_code_WB_reg_1_ ( .D(n5976), .CK(clk), .Q(
        pipeline_ctrl_prev_ex_code_WB[1]), .QN(n781) );
  DFF_X2 pipeline_ctrl_wfi_unkilled_WB_reg ( .D(n6207), .CK(clk), .QN(n9599)
         );
  DFF_X2 pipeline_ctrl_wr_reg_unkilled_WB_reg ( .D(n6252), .CK(clk), .Q(
        pipeline_ctrl_wr_reg_unkilled_WB), .QN(n791) );
  DFF_X2 pipeline_md_out_sel_reg_1_ ( .D(n6244), .CK(clk), .Q(
        pipeline_md_out_sel[1]), .QN(n1154) );
  DFF_X2 pipeline_md_op_reg_0_ ( .D(n6243), .CK(clk), .Q(pipeline_md_op_0_), 
        .QN(n963) );
  DFF_X2 pipeline_md_out_sel_reg_0_ ( .D(n6245), .CK(clk), .Q(
        pipeline_md_out_sel[0]), .QN(n1153) );
  DFF_X2 pipeline_md_b_reg_6_ ( .D(n5774), .CK(clk), .Q(pipeline_md_b[6]), 
        .QN(n12751) );
  DFF_X2 pipeline_md_result_reg_17_ ( .D(n5636), .CK(clk), .Q(
        pipeline_md_resp_result[17]) );
  DFF_X2 pipeline_md_result_reg_16_ ( .D(n5637), .CK(clk), .Q(
        pipeline_md_resp_result[16]) );
  DFF_X2 pipeline_md_result_reg_15_ ( .D(n5638), .CK(clk), .Q(
        pipeline_md_resp_result[15]) );
  DFF_X2 pipeline_md_result_reg_14_ ( .D(n5639), .CK(clk), .Q(
        pipeline_md_resp_result[14]) );
  DFF_X2 pipeline_md_result_reg_13_ ( .D(n5640), .CK(clk), .Q(
        pipeline_md_resp_result[13]) );
  DFF_X2 pipeline_md_result_reg_4_ ( .D(n5649), .CK(clk), .Q(
        pipeline_md_resp_result[4]) );
  DFF_X2 pipeline_md_result_reg_25_ ( .D(n5628), .CK(clk), .Q(
        pipeline_md_resp_result[25]) );
  DFF_X2 pipeline_md_result_reg_24_ ( .D(n5629), .CK(clk), .Q(
        pipeline_md_resp_result[24]) );
  DFF_X2 pipeline_md_result_reg_23_ ( .D(n5630), .CK(clk), .Q(
        pipeline_md_resp_result[23]) );
  DFF_X2 pipeline_md_result_reg_22_ ( .D(n5631), .CK(clk), .Q(
        pipeline_md_resp_result[22]) );
  DFF_X2 pipeline_md_result_reg_21_ ( .D(n5632), .CK(clk), .Q(
        pipeline_md_resp_result[21]) );
  DFF_X2 pipeline_md_result_reg_20_ ( .D(n5633), .CK(clk), .Q(
        pipeline_md_resp_result[20]) );
  DFF_X2 pipeline_md_result_reg_19_ ( .D(n5634), .CK(clk), .Q(
        pipeline_md_resp_result[19]) );
  DFF_X2 pipeline_md_result_reg_18_ ( .D(n5635), .CK(clk), .Q(
        pipeline_md_resp_result[18]) );
  DFF_X2 pipeline_md_result_reg_12_ ( .D(n5641), .CK(clk), .Q(
        pipeline_md_resp_result[12]) );
  DFF_X2 pipeline_md_result_reg_11_ ( .D(n5642), .CK(clk), .Q(
        pipeline_md_resp_result[11]) );
  DFF_X2 pipeline_md_result_reg_10_ ( .D(n5643), .CK(clk), .Q(
        pipeline_md_resp_result[10]) );
  DFF_X2 pipeline_md_result_reg_9_ ( .D(n5644), .CK(clk), .Q(
        pipeline_md_resp_result[9]) );
  DFF_X2 pipeline_md_result_reg_8_ ( .D(n5645), .CK(clk), .Q(
        pipeline_md_resp_result[8]) );
  DFF_X2 pipeline_md_result_reg_7_ ( .D(n5646), .CK(clk), .Q(
        pipeline_md_resp_result[7]) );
  DFF_X2 pipeline_md_result_reg_6_ ( .D(n5647), .CK(clk), .Q(
        pipeline_md_resp_result[6]) );
  DFF_X2 pipeline_md_result_reg_5_ ( .D(n5648), .CK(clk), .Q(
        pipeline_md_resp_result[5]) );
  DFF_X2 pipeline_md_result_reg_3_ ( .D(n5650), .CK(clk), .Q(
        pipeline_md_resp_result[3]) );
  DFF_X2 pipeline_md_result_reg_2_ ( .D(n5651), .CK(clk), .Q(
        pipeline_md_resp_result[2]) );
  DFF_X2 pipeline_md_result_reg_1_ ( .D(n5652), .CK(clk), .Q(
        pipeline_md_resp_result[1]) );
  DFF_X2 pipeline_md_result_reg_0_ ( .D(n5653), .CK(clk), .Q(
        pipeline_md_resp_result[0]) );
  DFF_X2 pipeline_csr_mtvec_reg_4_ ( .D(n6204), .CK(clk), .Q(
        pipeline_csr_mtvec[4]), .QN(n1195) );
  DFF_X2 pipeline_csr_mtvec_reg_3_ ( .D(n6205), .CK(clk), .Q(
        pipeline_csr_mtvec[3]), .QN(n10489) );
  DFF_X2 pipeline_alu_out_WB_reg_21_ ( .D(n5823), .CK(clk), .Q(
        pipeline_alu_out_WB[21]), .QN(n492) );
  DFF_X2 pipeline_alu_out_WB_reg_16_ ( .D(n5828), .CK(clk), .Q(
        pipeline_alu_out_WB[16]), .QN(n487) );
  DFF_X2 pipeline_csr_priv_stack_reg_4_ ( .D(n5981), .CK(clk), .QN(n12815) );
  DFF_X2 pipeline_csr_priv_stack_reg_3_ ( .D(n5982), .CK(clk), .QN(n12155) );
  DFF_X2 pipeline_csr_mtimecmp_reg_4_ ( .D(n6172), .CK(clk), .Q(
        pipeline_csr_mtimecmp[4]), .QN(n1291) );
  DFF_X2 pipeline_csr_from_host_reg_4_ ( .D(n6077), .CK(clk), .QN(n11234) );
  DFF_X2 pipeline_csr_mtvec_reg_6_ ( .D(n6202), .CK(clk), .Q(
        pipeline_csr_mtvec[6]), .QN(n1197) );
  DFF_X2 pipeline_csr_mie_reg_18_ ( .D(n6225), .CK(clk), .Q(
        pipeline_csr_mie[18]), .QN(n1533) );
  DFF_X2 pipeline_csr_mie_reg_13_ ( .D(n6220), .CK(clk), .Q(
        pipeline_csr_mie[13]), .QN(n1528) );
  DFF_X2 pipeline_csr_mie_reg_12_ ( .D(n6219), .CK(clk), .Q(
        pipeline_csr_mie[12]), .QN(n1527) );
  DFF_X2 pipeline_csr_mie_reg_11_ ( .D(n6218), .CK(clk), .Q(
        pipeline_csr_mie[11]), .QN(n1526) );
  DFF_X2 pipeline_csr_mie_reg_10_ ( .D(n6217), .CK(clk), .Q(
        pipeline_csr_mie[10]), .QN(n1525) );
  DFF_X2 pipeline_csr_to_host_reg_3_ ( .D(n6084), .CK(clk), .Q(
        pipeline_csr_to_host_3_), .QN(n1258) );
  DFF_X2 pipeline_csr_mtimecmp_reg_3_ ( .D(n6173), .CK(clk), .Q(
        pipeline_csr_mtimecmp[3]), .QN(n1290) );
  DFF_X2 pipeline_csr_from_host_reg_3_ ( .D(n6078), .CK(clk), .Q(
        pipeline_csr_from_host[3]), .QN(n1226) );
  DFF_X2 pipeline_alu_out_WB_reg_19_ ( .D(n5825), .CK(clk), .Q(
        pipeline_alu_out_WB[19]), .QN(n490) );
  DFF_X2 pipeline_alu_out_WB_reg_17_ ( .D(n5827), .CK(clk), .Q(
        pipeline_alu_out_WB[17]), .QN(n488) );
  DFF_X2 pipeline_csr_mtvec_reg_5_ ( .D(n6203), .CK(clk), .Q(
        pipeline_csr_mtvec[5]), .QN(n1196) );
  DFF_X2 pipeline_md_result_reg_26_ ( .D(n5627), .CK(clk), .Q(
        pipeline_md_resp_result[26]) );
  DFF_X2 pipeline_alu_out_WB_reg_20_ ( .D(n5824), .CK(clk), .Q(
        pipeline_alu_out_WB[20]), .QN(n491) );
  DFF_X2 pipeline_csr_from_host_reg_30_ ( .D(n6051), .CK(clk), .QN(n10249) );
  DFF_X2 pipeline_csr_from_host_reg_29_ ( .D(n6052), .CK(clk), .QN(n10365) );
  DFF_X2 pipeline_csr_from_host_reg_27_ ( .D(n6054), .CK(clk), .QN(n10468) );
  DFF_X2 pipeline_csr_from_host_reg_26_ ( .D(n6055), .CK(clk), .QN(n10544) );
  DFF_X2 pipeline_csr_from_host_reg_25_ ( .D(n6056), .CK(clk), .QN(n10598) );
  DFF_X2 pipeline_csr_from_host_reg_24_ ( .D(n6057), .CK(clk), .QN(n10652) );
  DFF_X2 pipeline_csr_from_host_reg_23_ ( .D(n6058), .CK(clk), .QN(n10706) );
  DFF_X2 pipeline_csr_from_host_reg_22_ ( .D(n6059), .CK(clk), .QN(n10757) );
  DFF_X2 pipeline_csr_from_host_reg_21_ ( .D(n6060), .CK(clk), .QN(n10842) );
  DFF_X2 pipeline_csr_from_host_reg_19_ ( .D(n6062), .CK(clk), .QN(n10950) );
  DFF_X2 pipeline_csr_from_host_reg_18_ ( .D(n6063), .CK(clk), .QN(n10997) );
  DFF_X2 pipeline_csr_from_host_reg_17_ ( .D(n6064), .CK(clk), .QN(n11057) );
  DFF_X2 pipeline_csr_from_host_reg_16_ ( .D(n6065), .CK(clk), .QN(n11084) );
  DFF_X2 pipeline_csr_from_host_reg_14_ ( .D(n6067), .CK(clk), .QN(n11142) );
  DFF_X2 pipeline_csr_from_host_reg_13_ ( .D(n6068), .CK(clk), .QN(n11030) );
  DFF_X2 pipeline_csr_from_host_reg_12_ ( .D(n6069), .CK(clk), .QN(n10869) );
  DFF_X2 pipeline_csr_from_host_reg_11_ ( .D(n6070), .CK(clk), .QN(n10923) );
  DFF_X2 pipeline_csr_from_host_reg_10_ ( .D(n6071), .CK(clk), .QN(n10977) );
  DFF_X2 pipeline_csr_from_host_reg_9_ ( .D(n6072), .CK(clk), .QN(n10571) );
  DFF_X2 pipeline_csr_mtimecmp_reg_30_ ( .D(n6146), .CK(clk), .Q(
        pipeline_csr_mtimecmp[30]), .QN(n10243) );
  DFF_X2 pipeline_csr_mtimecmp_reg_29_ ( .D(n6147), .CK(clk), .Q(
        pipeline_csr_mtimecmp[29]), .QN(n10362) );
  DFF_X2 pipeline_csr_mtimecmp_reg_27_ ( .D(n6149), .CK(clk), .Q(
        pipeline_csr_mtimecmp[27]), .QN(n10465) );
  DFF_X2 pipeline_csr_mtimecmp_reg_26_ ( .D(n6150), .CK(clk), .Q(
        pipeline_csr_mtimecmp[26]), .QN(n10541) );
  DFF_X2 pipeline_csr_mtimecmp_reg_25_ ( .D(n6151), .CK(clk), .Q(
        pipeline_csr_mtimecmp[25]), .QN(n10595) );
  DFF_X2 pipeline_csr_mtimecmp_reg_24_ ( .D(n6152), .CK(clk), .Q(
        pipeline_csr_mtimecmp[24]), .QN(n10649) );
  DFF_X2 pipeline_csr_mtimecmp_reg_23_ ( .D(n6153), .CK(clk), .Q(
        pipeline_csr_mtimecmp[23]), .QN(n10703) );
  DFF_X2 pipeline_csr_mtimecmp_reg_22_ ( .D(n6154), .CK(clk), .Q(
        pipeline_csr_mtimecmp[22]), .QN(n10754) );
  DFF_X2 pipeline_csr_mtimecmp_reg_21_ ( .D(n6155), .CK(clk), .Q(
        pipeline_csr_mtimecmp[21]), .QN(n10839) );
  DFF_X2 pipeline_csr_mtimecmp_reg_20_ ( .D(n6156), .CK(clk), .Q(
        pipeline_csr_mtimecmp[20]), .QN(n10891) );
  DFF_X2 pipeline_csr_mtimecmp_reg_19_ ( .D(n6157), .CK(clk), .Q(
        pipeline_csr_mtimecmp[19]), .QN(n10947) );
  DFF_X2 pipeline_csr_mtimecmp_reg_18_ ( .D(n6158), .CK(clk), .Q(
        pipeline_csr_mtimecmp[18]), .QN(n11005) );
  DFF_X2 pipeline_csr_mtimecmp_reg_17_ ( .D(n6159), .CK(clk), .Q(
        pipeline_csr_mtimecmp[17]), .QN(n11054) );
  DFF_X2 pipeline_csr_mtimecmp_reg_16_ ( .D(n6160), .CK(clk), .Q(
        pipeline_csr_mtimecmp[16]), .QN(n11081) );
  DFF_X2 pipeline_csr_mtimecmp_reg_15_ ( .D(n6161), .CK(clk), .Q(
        pipeline_csr_mtimecmp[15]), .QN(n11107) );
  DFF_X2 pipeline_csr_mtimecmp_reg_14_ ( .D(n6162), .CK(clk), .Q(
        pipeline_csr_mtimecmp[14]), .QN(n11139) );
  DFF_X2 pipeline_csr_mtimecmp_reg_13_ ( .D(n6163), .CK(clk), .Q(
        pipeline_csr_mtimecmp[13]), .QN(n11027) );
  DFF_X2 pipeline_csr_mtimecmp_reg_12_ ( .D(n6164), .CK(clk), .Q(
        pipeline_csr_mtimecmp[12]), .QN(n10866) );
  DFF_X2 pipeline_csr_mtimecmp_reg_11_ ( .D(n6165), .CK(clk), .Q(
        pipeline_csr_mtimecmp[11]), .QN(n10920) );
  DFF_X2 pipeline_csr_mtimecmp_reg_10_ ( .D(n6166), .CK(clk), .Q(
        pipeline_csr_mtimecmp[10]), .QN(n10974) );
  DFF_X2 pipeline_csr_mtimecmp_reg_9_ ( .D(n6167), .CK(clk), .Q(
        pipeline_csr_mtimecmp[9]), .QN(n10568) );
  DFF_X2 pipeline_csr_mtimecmp_reg_6_ ( .D(n6170), .CK(clk), .Q(
        pipeline_csr_mtimecmp[6]), .QN(n10731) );
  DFF_X2 pipeline_csr_mscratch_reg_30_ ( .D(n6114), .CK(clk), .Q(
        pipeline_csr_mscratch[30]), .QN(n1191) );
  DFF_X2 pipeline_csr_mscratch_reg_29_ ( .D(n6115), .CK(clk), .Q(
        pipeline_csr_mscratch[29]), .QN(n1190) );
  DFF_X2 pipeline_csr_mscratch_reg_27_ ( .D(n6117), .CK(clk), .Q(
        pipeline_csr_mscratch[27]), .QN(n1188) );
  DFF_X2 pipeline_csr_mscratch_reg_26_ ( .D(n6118), .CK(clk), .Q(
        pipeline_csr_mscratch[26]), .QN(n1187) );
  DFF_X2 pipeline_csr_mscratch_reg_25_ ( .D(n6119), .CK(clk), .Q(
        pipeline_csr_mscratch[25]), .QN(n1186) );
  DFF_X2 pipeline_csr_mscratch_reg_24_ ( .D(n6120), .CK(clk), .Q(
        pipeline_csr_mscratch[24]), .QN(n1185) );
  DFF_X2 pipeline_csr_mscratch_reg_23_ ( .D(n6121), .CK(clk), .Q(
        pipeline_csr_mscratch[23]), .QN(n1184) );
  DFF_X2 pipeline_csr_mscratch_reg_22_ ( .D(n6122), .CK(clk), .Q(
        pipeline_csr_mscratch[22]), .QN(n1183) );
  DFF_X2 pipeline_csr_mscratch_reg_21_ ( .D(n6123), .CK(clk), .Q(
        pipeline_csr_mscratch[21]), .QN(n1182) );
  DFF_X2 pipeline_csr_mscratch_reg_20_ ( .D(n6124), .CK(clk), .Q(
        pipeline_csr_mscratch[20]), .QN(n1181) );
  DFF_X2 pipeline_csr_mscratch_reg_19_ ( .D(n6125), .CK(clk), .Q(
        pipeline_csr_mscratch[19]), .QN(n1180) );
  DFF_X2 pipeline_csr_mscratch_reg_18_ ( .D(n6126), .CK(clk), .Q(
        pipeline_csr_mscratch[18]), .QN(n1179) );
  DFF_X2 pipeline_csr_mscratch_reg_17_ ( .D(n6127), .CK(clk), .Q(
        pipeline_csr_mscratch[17]), .QN(n1178) );
  DFF_X2 pipeline_csr_mscratch_reg_16_ ( .D(n6128), .CK(clk), .Q(
        pipeline_csr_mscratch[16]), .QN(n1177) );
  DFF_X2 pipeline_csr_mscratch_reg_15_ ( .D(n6129), .CK(clk), .Q(
        pipeline_csr_mscratch[15]), .QN(n1176) );
  DFF_X2 pipeline_csr_mscratch_reg_14_ ( .D(n6130), .CK(clk), .Q(
        pipeline_csr_mscratch[14]), .QN(n1175) );
  DFF_X2 pipeline_csr_mscratch_reg_13_ ( .D(n6131), .CK(clk), .Q(
        pipeline_csr_mscratch[13]), .QN(n1174) );
  DFF_X2 pipeline_csr_mscratch_reg_12_ ( .D(n6132), .CK(clk), .Q(
        pipeline_csr_mscratch[12]), .QN(n1173) );
  DFF_X2 pipeline_csr_mscratch_reg_11_ ( .D(n6133), .CK(clk), .Q(
        pipeline_csr_mscratch[11]), .QN(n1172) );
  DFF_X2 pipeline_csr_mscratch_reg_10_ ( .D(n6134), .CK(clk), .Q(
        pipeline_csr_mscratch[10]), .QN(n1171) );
  DFF_X2 pipeline_csr_mscratch_reg_9_ ( .D(n6135), .CK(clk), .Q(
        pipeline_csr_mscratch[9]), .QN(n1170) );
  DFF_X2 pipeline_csr_mscratch_reg_6_ ( .D(n6138), .CK(clk), .Q(
        pipeline_csr_mscratch[6]), .QN(n1167) );
  DFF_X2 pipeline_csr_from_host_reg_28_ ( .D(n6053), .CK(clk), .Q(
        pipeline_csr_from_host[28]), .QN(n1251) );
  DFF_X2 pipeline_csr_mtimecmp_reg_28_ ( .D(n6148), .CK(clk), .Q(
        pipeline_csr_mtimecmp[28]), .QN(n10430) );
  DFF_X2 pipeline_csr_mscratch_reg_28_ ( .D(n6116), .CK(clk), .Q(
        pipeline_csr_mscratch[28]), .QN(n1189) );
  DFF_X2 pipeline_csr_priv_stack_reg_5_ ( .D(n5980), .CK(clk), .QN(n12821) );
  DFF_X2 pipeline_csr_mtimecmp_reg_5_ ( .D(n6171), .CK(clk), .Q(
        pipeline_csr_mtimecmp[5]), .QN(n1292) );
  DFF_X2 pipeline_csr_from_host_reg_5_ ( .D(n6076), .CK(clk), .Q(
        pipeline_csr_from_host[5]), .QN(n1228) );
  DFF_X2 pipeline_alu_out_WB_reg_18_ ( .D(n5826), .CK(clk), .Q(
        pipeline_alu_out_WB[18]), .QN(n489) );
  DFF_X2 pipeline_alu_out_WB_reg_14_ ( .D(n5830), .CK(clk), .Q(
        pipeline_alu_out_WB[14]), .QN(n485) );
  DFF_X2 pipeline_csr_instret_full_reg_36_ ( .D(n6010), .CK(clk), .Q(
        pipeline_csr_instret_full[36]), .QN(n11231) );
  DFF_X2 pipeline_csr_instret_full_reg_4_ ( .D(n6042), .CK(clk), .Q(
        pipeline_csr_instret_full[4]), .QN(n1387) );
  DFF_X2 pipeline_csr_instret_full_reg_35_ ( .D(n6011), .CK(clk), .Q(
        pipeline_csr_instret_full[35]), .QN(n1418) );
  DFF_X2 pipeline_csr_instret_full_reg_3_ ( .D(n6043), .CK(clk), .Q(
        pipeline_csr_instret_full[3]), .QN(n10492) );
  DFF_X2 pipeline_csr_mbadaddr_reg_16_ ( .D(n5796), .CK(clk), .QN(n11382) );
  DFF_X2 pipeline_csr_mbadaddr_reg_15_ ( .D(n5797), .CK(clk), .QN(n11352) );
  DFF_X2 pipeline_csr_mbadaddr_reg_14_ ( .D(n5798), .CK(clk), .QN(n11194) );
  DFF_X2 pipeline_csr_mbadaddr_reg_17_ ( .D(n5795), .CK(clk), .QN(n11421) );
  DFF_X2 pipeline_csr_mtvec_reg_2_ ( .D(n6206), .CK(clk), .Q(
        pipeline_csr_mtvec[2]), .QN(n1193) );
  DFF_X2 pipeline_csr_mbadaddr_reg_22_ ( .D(n5790), .CK(clk), .QN(n11785) );
  DFF_X2 pipeline_csr_mbadaddr_reg_18_ ( .D(n5794), .CK(clk), .QN(n11481) );
  DFF_X2 pipeline_csr_mbadaddr_reg_21_ ( .D(n5791), .CK(clk), .QN(n11701) );
  DFF_X2 pipeline_csr_mbadaddr_reg_20_ ( .D(n5792), .CK(clk), .QN(n11627) );
  DFF_X2 pipeline_csr_mbadaddr_reg_13_ ( .D(n5799), .CK(clk), .QN(n11451) );
  DFF_X2 pipeline_csr_mbadaddr_reg_23_ ( .D(n5789), .CK(clk), .QN(n11855) );
  DFF_X2 pipeline_csr_mbadaddr_reg_5_ ( .D(n5807), .CK(clk), .QN(n11737) );
  DFF_X2 pipeline_alu_out_WB_reg_7_ ( .D(n5837), .CK(clk), .Q(
        pipeline_alu_out_WB[7]), .QN(n478) );
  DFF_X2 pipeline_csr_from_host_reg_31_ ( .D(n6050), .CK(clk), .Q(
        pipeline_csr_from_host[31]), .QN(n1254) );
  DFF_X2 pipeline_csr_mtimecmp_reg_31_ ( .D(n6145), .CK(clk), .Q(
        pipeline_csr_mtimecmp[31]), .QN(n10287) );
  DFF_X2 pipeline_csr_mscratch_reg_31_ ( .D(n6113), .CK(clk), .Q(
        pipeline_csr_mscratch[31]), .QN(n1192) );
  DFF_X2 pipeline_csr_mbadaddr_reg_6_ ( .D(n5806), .CK(clk), .QN(n11814) );
  DFF_X2 pipeline_csr_mbadaddr_reg_11_ ( .D(n5801), .CK(clk), .QN(n11593) );
  DFF_X2 pipeline_csr_mbadaddr_reg_29_ ( .D(n5783), .CK(clk), .QN(n12328) );
  DFF_X2 pipeline_csr_mbadaddr_reg_28_ ( .D(n5784), .CK(clk), .QN(n12232) );
  DFF_X2 pipeline_csr_mie_reg_8_ ( .D(n6215), .CK(clk), .Q(pipeline_csr_mie[8]), .QN(n1523) );
  DFF_X2 pipeline_csr_mbadaddr_reg_19_ ( .D(n5793), .CK(clk), .QN(n11555) );
  DFF_X2 pipeline_csr_mbadaddr_reg_10_ ( .D(n5802), .CK(clk), .QN(n11517) );
  DFF_X2 pipeline_csr_mbadaddr_reg_25_ ( .D(n5787), .CK(clk), .QN(n12040) );
  DFF_X2 pipeline_csr_mbadaddr_reg_24_ ( .D(n5788), .CK(clk), .QN(n11970) );
  DFF_X2 pipeline_csr_mbadaddr_reg_26_ ( .D(n5786), .CK(clk), .QN(n12108) );
  DFF_X2 pipeline_csr_mbadaddr_reg_9_ ( .D(n5803), .CK(clk), .QN(n12072) );
  DFF_X2 pipeline_csr_mbadaddr_reg_12_ ( .D(n5800), .CK(clk), .QN(n11660) );
  DFF_X2 pipeline_csr_mbadaddr_reg_30_ ( .D(n5782), .CK(clk), .QN(n12665) );
  DFF_X2 pipeline_csr_mbadaddr_reg_0_ ( .D(n5812), .CK(clk), .Q(
        pipeline_csr_mbadaddr[0]), .QN(n1447) );
  DFF_X2 pipeline_csr_mie_reg_7_ ( .D(n6214), .CK(clk), .Q(pipeline_csr_mie[7]), .QN(n1522) );
  DFF_X2 pipeline_csr_mbadaddr_reg_27_ ( .D(n5785), .CK(clk), .QN(n12186) );
  DFF_X2 pipeline_alu_out_WB_reg_22_ ( .D(n5822), .CK(clk), .Q(
        pipeline_alu_out_WB[22]), .QN(n493) );
  DFF_X2 pipeline_csr_priv_stack_reg_2_ ( .D(n6296), .CK(clk), .Q(
        pipeline_ctrl_N82), .QN(n10407) );
  DFF_X2 pipeline_alu_out_WB_reg_11_ ( .D(n5833), .CK(clk), .Q(
        pipeline_alu_out_WB[11]), .QN(n482) );
  DFF_X2 pipeline_csr_instret_full_reg_30_ ( .D(n6016), .CK(clk), .Q(
        pipeline_csr_instret_full[30]), .QN(n10252) );
  DFF_X2 pipeline_csr_instret_full_reg_29_ ( .D(n6017), .CK(clk), .Q(
        pipeline_csr_instret_full[29]), .QN(n10367) );
  DFF_X2 pipeline_csr_instret_full_reg_58_ ( .D(n5988), .CK(clk), .Q(
        pipeline_csr_instret_full[58]), .QN(n1441) );
  DFF_X2 pipeline_csr_instret_full_reg_57_ ( .D(n5989), .CK(clk), .Q(
        pipeline_csr_instret_full[57]), .QN(n1440) );
  DFF_X2 pipeline_csr_instret_full_reg_56_ ( .D(n5990), .CK(clk), .Q(
        pipeline_csr_instret_full[56]), .QN(n1439) );
  DFF_X2 pipeline_csr_instret_full_reg_55_ ( .D(n5991), .CK(clk), .Q(
        pipeline_csr_instret_full[55]), .QN(n1438) );
  DFF_X2 pipeline_csr_instret_full_reg_54_ ( .D(n5992), .CK(clk), .Q(
        pipeline_csr_instret_full[54]), .QN(n10758) );
  DFF_X2 pipeline_csr_instret_full_reg_53_ ( .D(n5993), .CK(clk), .Q(
        pipeline_csr_instret_full[53]), .QN(n10843) );
  DFF_X2 pipeline_csr_instret_full_reg_51_ ( .D(n5995), .CK(clk), .Q(
        pipeline_csr_instret_full[51]), .QN(n10951) );
  DFF_X2 pipeline_csr_instret_full_reg_50_ ( .D(n5996), .CK(clk), .Q(
        pipeline_csr_instret_full[50]), .QN(n10998) );
  DFF_X2 pipeline_csr_instret_full_reg_49_ ( .D(n5997), .CK(clk), .Q(
        pipeline_csr_instret_full[49]), .QN(n11058) );
  DFF_X2 pipeline_csr_instret_full_reg_48_ ( .D(n5998), .CK(clk), .Q(
        pipeline_csr_instret_full[48]), .QN(n11085) );
  DFF_X2 pipeline_csr_instret_full_reg_46_ ( .D(n6000), .CK(clk), .Q(
        pipeline_csr_instret_full[46]), .QN(n11143) );
  DFF_X2 pipeline_csr_instret_full_reg_45_ ( .D(n6001), .CK(clk), .Q(
        pipeline_csr_instret_full[45]), .QN(n11031) );
  DFF_X2 pipeline_csr_instret_full_reg_44_ ( .D(n6002), .CK(clk), .Q(
        pipeline_csr_instret_full[44]), .QN(n10870) );
  DFF_X2 pipeline_csr_instret_full_reg_43_ ( .D(n6003), .CK(clk), .Q(
        pipeline_csr_instret_full[43]), .QN(n10924) );
  DFF_X2 pipeline_csr_instret_full_reg_42_ ( .D(n6004), .CK(clk), .Q(
        pipeline_csr_instret_full[42]), .QN(n10978) );
  DFF_X2 pipeline_csr_instret_full_reg_41_ ( .D(n6005), .CK(clk), .Q(
        pipeline_csr_instret_full[41]), .QN(n10572) );
  DFF_X2 pipeline_csr_instret_full_reg_38_ ( .D(n6008), .CK(clk), .Q(
        pipeline_csr_instret_full[38]), .QN(n10733) );
  DFF_X2 pipeline_csr_instret_full_reg_27_ ( .D(n6019), .CK(clk), .Q(
        pipeline_csr_instret_full[27]), .QN(n10470) );
  DFF_X2 pipeline_csr_instret_full_reg_26_ ( .D(n6020), .CK(clk), .Q(
        pipeline_csr_instret_full[26]), .QN(n10546) );
  DFF_X2 pipeline_csr_instret_full_reg_25_ ( .D(n6021), .CK(clk), .Q(
        pipeline_csr_instret_full[25]), .QN(n10600) );
  DFF_X2 pipeline_csr_instret_full_reg_24_ ( .D(n6022), .CK(clk), .Q(
        pipeline_csr_instret_full[24]), .QN(n10654) );
  DFF_X2 pipeline_csr_instret_full_reg_23_ ( .D(n6023), .CK(clk), .Q(
        pipeline_csr_instret_full[23]), .QN(n10708) );
  DFF_X2 pipeline_csr_instret_full_reg_22_ ( .D(n6024), .CK(clk), .Q(
        pipeline_csr_instret_full[22]), .QN(n10760) );
  DFF_X2 pipeline_csr_instret_full_reg_21_ ( .D(n6025), .CK(clk), .Q(
        pipeline_csr_instret_full[21]), .QN(n10845) );
  DFF_X2 pipeline_csr_instret_full_reg_20_ ( .D(n6026), .CK(clk), .Q(
        pipeline_csr_instret_full[20]), .QN(n10893) );
  DFF_X2 pipeline_csr_instret_full_reg_19_ ( .D(n6027), .CK(clk), .Q(
        pipeline_csr_instret_full[19]), .QN(n10953) );
  DFF_X2 pipeline_csr_instret_full_reg_18_ ( .D(n6028), .CK(clk), .Q(
        pipeline_csr_instret_full[18]), .QN(n11000) );
  DFF_X2 pipeline_csr_instret_full_reg_17_ ( .D(n6029), .CK(clk), .Q(
        pipeline_csr_instret_full[17]), .QN(n11060) );
  DFF_X2 pipeline_csr_instret_full_reg_16_ ( .D(n6030), .CK(clk), .Q(
        pipeline_csr_instret_full[16]), .QN(n11087) );
  DFF_X2 pipeline_csr_instret_full_reg_15_ ( .D(n6031), .CK(clk), .Q(
        pipeline_csr_instret_full[15]), .QN(n11109) );
  DFF_X2 pipeline_csr_instret_full_reg_14_ ( .D(n6032), .CK(clk), .Q(
        pipeline_csr_instret_full[14]), .QN(n11145) );
  DFF_X2 pipeline_csr_instret_full_reg_13_ ( .D(n6033), .CK(clk), .Q(
        pipeline_csr_instret_full[13]), .QN(n11033) );
  DFF_X2 pipeline_csr_instret_full_reg_12_ ( .D(n6034), .CK(clk), .Q(
        pipeline_csr_instret_full[12]), .QN(n10872) );
  DFF_X2 pipeline_csr_instret_full_reg_11_ ( .D(n6035), .CK(clk), .Q(
        pipeline_csr_instret_full[11]), .QN(n10926) );
  DFF_X2 pipeline_csr_instret_full_reg_10_ ( .D(n6036), .CK(clk), .Q(
        pipeline_csr_instret_full[10]), .QN(n10980) );
  DFF_X2 pipeline_csr_instret_full_reg_9_ ( .D(n6037), .CK(clk), .Q(
        pipeline_csr_instret_full[9]), .QN(n10574) );
  DFF_X2 pipeline_csr_instret_full_reg_61_ ( .D(n6047), .CK(clk), .Q(
        pipeline_csr_instret_full[61]), .QN(n1444) );
  DFF_X2 pipeline_csr_instret_full_reg_59_ ( .D(n5987), .CK(clk), .Q(
        pipeline_csr_instret_full[59]), .QN(n1442) );
  DFF_X2 pipeline_csr_instret_full_reg_28_ ( .D(n6018), .CK(clk), .Q(
        pipeline_csr_instret_full[28]), .QN(n10433) );
  DFF_X2 pipeline_csr_instret_full_reg_60_ ( .D(n5986), .CK(clk), .Q(
        pipeline_csr_instret_full[60]), .QN(n1443) );
  DFF_X2 pipeline_md_result_reg_27_ ( .D(n5626), .CK(clk), .Q(
        pipeline_md_resp_result[27]) );
  DFF_X2 pipeline_csr_instret_full_reg_37_ ( .D(n6009), .CK(clk), .Q(
        pipeline_csr_instret_full[37]), .QN(n1420) );
  DFF_X2 pipeline_csr_instret_full_reg_5_ ( .D(n6041), .CK(clk), .Q(
        pipeline_csr_instret_full[5]), .QN(n10785) );
  DFF_X2 pipeline_csr_mbadaddr_reg_7_ ( .D(n5805), .CK(clk), .QN(n11890) );
  DFF_X2 pipeline_csr_mie_reg_31_ ( .D(n6238), .CK(clk), .Q(
        pipeline_csr_mie[31]), .QN(n1546) );
  DFF_X2 pipeline_csr_mtimecmp_reg_8_ ( .D(n6168), .CK(clk), .Q(
        pipeline_csr_mtimecmp[8]), .QN(n10620) );
  DFF_X2 pipeline_csr_mscratch_reg_8_ ( .D(n6136), .CK(clk), .Q(
        pipeline_csr_mscratch[8]), .QN(n1169) );
  DFF_X2 pipeline_csr_mbadaddr_reg_4_ ( .D(n5808), .CK(clk), .QN(n12804) );
  DFF_X2 pipeline_csr_from_host_reg_7_ ( .D(n6074), .CK(clk), .QN(n10680) );
  DFF_X2 pipeline_csr_mtimecmp_reg_7_ ( .D(n6169), .CK(clk), .Q(
        pipeline_csr_mtimecmp[7]), .QN(n10677) );
  DFF_X2 pipeline_csr_mscratch_reg_7_ ( .D(n6137), .CK(clk), .Q(
        pipeline_csr_mscratch[7]), .QN(n1168) );
  DFF_X2 pipeline_alu_out_WB_reg_23_ ( .D(n5821), .CK(clk), .Q(
        pipeline_alu_out_WB[23]), .QN(n494) );
  DFF_X2 pipeline_csr_mbadaddr_reg_8_ ( .D(n5804), .CK(clk), .QN(n11997) );
  DFF_X2 pipeline_csr_mtimecmp_reg_2_ ( .D(n6174), .CK(clk), .Q(
        pipeline_csr_mtimecmp[2]), .QN(n1289) );
  DFF_X2 pipeline_csr_from_host_reg_2_ ( .D(n6079), .CK(clk), .QN(n10401) );
  DFF_X2 pipeline_csr_instret_full_reg_62_ ( .D(n5985), .CK(clk), .Q(
        pipeline_csr_instret_full[62]), .QN(n1445) );
  DFF_X2 pipeline_csr_instret_full_reg_0_ ( .D(n6046), .CK(clk), .Q(
        pipeline_csr_instret_full[0]), .QN(n1319) );
  DFF_X2 pipeline_csr_priv_stack_reg_0_ ( .D(n6297), .CK(clk), .Q(
        pipeline_csr_priv_stack_0), .QN(n1549) );
  DFF_X2 pipeline_csr_msip_reg ( .D(n6240), .CK(clk), .Q(pipeline_csr_mip_3), 
        .QN(n10510) );
  DFF_X2 pipeline_csr_instret_full_reg_31_ ( .D(n6015), .CK(clk), .Q(
        pipeline_csr_instret_full[31]), .QN(n10293) );
  DFF_X2 pipeline_csr_mtimecmp_reg_0_ ( .D(n6176), .CK(clk), .Q(
        pipeline_csr_mtimecmp[0]), .QN(n1287) );
  DFF_X2 pipeline_csr_from_host_reg_0_ ( .D(n6081), .CK(clk), .Q(
        pipeline_csr_from_host[0]), .QN(n1223) );
  DFF_X2 pipeline_csr_instret_full_reg_34_ ( .D(n6012), .CK(clk), .Q(
        pipeline_csr_instret_full[34]), .QN(n10399) );
  DFF_X2 pipeline_csr_instret_full_reg_2_ ( .D(n6044), .CK(clk), .Q(
        pipeline_csr_instret_full[2]), .QN(n1385) );
  DFF_X2 pipeline_alu_out_WB_reg_15_ ( .D(n5829), .CK(clk), .Q(
        pipeline_alu_out_WB[15]), .QN(n486) );
  DFF_X2 pipeline_csr_instret_full_reg_8_ ( .D(n6038), .CK(clk), .Q(
        pipeline_csr_instret_full[8]), .QN(n10622) );
  DFF_X2 pipeline_csr_instret_full_reg_39_ ( .D(n6007), .CK(clk), .Q(
        pipeline_csr_instret_full[39]), .QN(n1422) );
  DFF_X2 pipeline_csr_instret_full_reg_7_ ( .D(n6039), .CK(clk), .Q(
        pipeline_csr_instret_full[7]), .QN(n10682) );
  DFF_X2 pipeline_md_result_reg_28_ ( .D(n5625), .CK(clk), .Q(
        pipeline_md_resp_result[28]) );
  DFF_X2 pipeline_csr_instret_full_reg_63_ ( .D(n5984), .CK(clk), .Q(
        pipeline_csr_instret_full[63]), .QN(n10292) );
  DFF_X2 pipeline_csr_mbadaddr_reg_31_ ( .D(n5781), .CK(clk), .QN(n12595) );
  DFF_X2 pipeline_alu_out_WB_reg_12_ ( .D(n5832), .CK(clk), .Q(
        pipeline_alu_out_WB[12]), .QN(n483) );
  DFF_X2 pipeline_csr_instret_full_reg_32_ ( .D(n6014), .CK(clk), .Q(
        pipeline_csr_instret_full[32]), .QN(n11259) );
  DFF_X2 pipeline_alu_out_WB_reg_3_ ( .D(n5841), .CK(clk), .Q(
        pipeline_alu_out_WB[3]), .QN(n474) );
  DFF_X2 pipeline_alu_out_WB_reg_25_ ( .D(n5819), .CK(clk), .Q(
        pipeline_alu_out_WB[25]), .QN(n496) );
  DFF_X2 pipeline_csr_mbadaddr_reg_2_ ( .D(n5810), .CK(clk), .QN(n12288) );
  DFF_X2 pipeline_alu_out_WB_reg_13_ ( .D(n5831), .CK(clk), .Q(
        pipeline_alu_out_WB[13]), .QN(n484) );
  DFF_X2 pipeline_alu_out_WB_reg_0_ ( .D(n6301), .CK(clk), .Q(
        pipeline_alu_out_WB[0]), .QN(n12937) );
  DFF_X2 pipeline_ctrl_had_ex_DX_reg ( .D(n6300), .CK(clk), .Q(
        pipeline_ctrl_had_ex_DX), .QN(n799) );
  DFF_X2 pipeline_alu_out_WB_reg_4_ ( .D(n5840), .CK(clk), .Q(
        pipeline_alu_out_WB[4]), .QN(n475) );
  DFF_X2 pipeline_alu_out_WB_reg_8_ ( .D(n5836), .CK(clk), .Q(
        pipeline_alu_out_WB[8]), .QN(n479) );
  DFF_X2 pipeline_alu_out_WB_reg_10_ ( .D(n5834), .CK(clk), .Q(
        pipeline_alu_out_WB[10]), .QN(n481) );
  DFF_X2 pipeline_md_result_reg_29_ ( .D(n5624), .CK(clk), .Q(
        pipeline_md_resp_result[29]) );
  DFF_X2 pipeline_alu_out_WB_reg_9_ ( .D(n5835), .CK(clk), .Q(
        pipeline_alu_out_WB[9]), .QN(n480) );
  DFF_X2 pipeline_alu_out_WB_reg_5_ ( .D(n5839), .CK(clk), .Q(
        pipeline_alu_out_WB[5]), .QN(n476) );
  DFF_X2 pipeline_alu_out_WB_reg_6_ ( .D(n5838), .CK(clk), .Q(
        pipeline_alu_out_WB[6]), .QN(n477) );
  DFF_X2 pipeline_alu_out_WB_reg_24_ ( .D(n5820), .CK(clk), .Q(
        pipeline_alu_out_WB[24]), .QN(n495) );
  DFF_X2 pipeline_csr_priv_stack_reg_1_ ( .D(n6298), .CK(clk), .Q(
        pipeline_ctrl_N81), .QN(n10323) );
  DFF_X2 pipeline_csr_instret_full_reg_33_ ( .D(n6013), .CK(clk), .Q(
        pipeline_csr_instret_full[33]), .QN(n10317) );
  DFF_X2 pipeline_csr_instret_full_reg_1_ ( .D(n6045), .CK(clk), .Q(
        pipeline_csr_instret_full[1]), .QN(n1384) );
  DFF_X2 pipeline_md_result_reg_30_ ( .D(n5623), .CK(clk), .Q(
        pipeline_md_resp_result[30]) );
  DFF_X2 pipeline_csr_mtip_reg ( .D(n6366), .CK(clk), .Q(pipeline_csr_mip_7_), 
        .QN(n1547) );
  DFF_X2 pipeline_csr_mtimecmp_reg_1_ ( .D(n6175), .CK(clk), .Q(
        pipeline_csr_mtimecmp[1]), .QN(n1288) );
  DFF_X2 pipeline_csr_from_host_reg_1_ ( .D(n6080), .CK(clk), .Q(
        pipeline_csr_from_host[1]), .QN(n1224) );
  DFF_X2 pipeline_alu_out_WB_reg_2_ ( .D(n5842), .CK(clk), .Q(
        pipeline_alu_out_WB[2]), .QN(n473) );
  DFF_X2 pipeline_alu_out_WB_reg_26_ ( .D(n5818), .CK(clk), .Q(
        pipeline_alu_out_WB[26]), .QN(n497) );
  DFF_X2 pipeline_csr_mbadaddr_reg_1_ ( .D(n5811), .CK(clk), .Q(
        pipeline_csr_mbadaddr[1]), .QN(n1448) );
  DFF_X2 pipeline_md_result_reg_31_ ( .D(n5622), .CK(clk), .Q(
        pipeline_md_resp_result[31]) );
  DFF_X2 pipeline_alu_out_WB_reg_1_ ( .D(n5843), .CK(clk), .Q(
        pipeline_alu_out_WB[1]), .QN(n12936) );
  DFF_X2 pipeline_ctrl_prev_killed_DX_reg ( .D(n6049), .CK(clk), .Q(
        pipeline_ctrl_prev_killed_DX), .QN(n800) );
  DFF_X2 pipeline_inst_DX_reg_4_ ( .D(n6259), .CK(clk), .Q(pipeline_inst_DX[4]), .QN(n9631) );
  DFF_X2 pipeline_alu_out_WB_reg_27_ ( .D(n5817), .CK(clk), .Q(
        pipeline_alu_out_WB[27]), .QN(n498) );
  DFF_X2 pipeline_inst_DX_reg_23_ ( .D(n6286), .CK(clk), .Q(
        pipeline_regfile_N20), .QN(n8223) );
  DFF_X2 pipeline_inst_DX_reg_28_ ( .D(n6291), .CK(clk), .Q(
        pipeline_inst_DX[28]), .QN(n9634) );
  DFF_X2 pipeline_inst_DX_reg_29_ ( .D(n6292), .CK(clk), .Q(
        pipeline_inst_DX[29]), .QN(n9632) );
  DFF_X2 pipeline_PC_IF_reg_1_ ( .D(n5970), .CK(clk), .QN(n12535) );
  DFF_X2 pipeline_inst_DX_reg_3_ ( .D(n6258), .CK(clk), .Q(pipeline_inst_DX[3]), .QN(n9648) );
  DFF_X2 pipeline_inst_DX_reg_25_ ( .D(n6288), .CK(clk), .Q(
        pipeline_inst_DX[25]), .QN(n10336) );
  DFF_X2 pipeline_inst_DX_reg_31_ ( .D(n6295), .CK(clk), .Q(pipeline_imm_31_), 
        .QN(n10242) );
  DFF_X2 pipeline_inst_DX_reg_6_ ( .D(n6261), .CK(clk), .Q(pipeline_inst_DX[6]), .QN(n9650) );
  DFF_X2 pipeline_inst_DX_reg_24_ ( .D(n6287), .CK(clk), .Q(
        pipeline_regfile_N21), .QN(n8214) );
  DFF_X2 pipeline_inst_DX_reg_5_ ( .D(n6260), .CK(clk), .Q(pipeline_inst_DX[5]), .QN(n9651) );
  DFF_X2 pipeline_inst_DX_reg_2_ ( .D(n6257), .CK(clk), .Q(pipeline_inst_DX[2]), .QN(n9623) );
  DFF_X2 pipeline_inst_DX_reg_26_ ( .D(n6289), .CK(clk), .Q(n10235), .QN(
        n10338) );
  DFF_X2 pipeline_inst_DX_reg_19_ ( .D(n6282), .CK(clk), .Q(
        pipeline_regfile_N16), .QN(n9270) );
  DFF_X2 pipeline_inst_DX_reg_18_ ( .D(n6281), .CK(clk), .Q(
        pipeline_regfile_N15), .QN(n9279) );
  DFF_X2 pipeline_inst_DX_reg_27_ ( .D(n6290), .CK(clk), .Q(n10337), .QN(
        n10236) );
  DFF_X2 pipeline_PC_DX_reg_30_ ( .D(n5879), .CK(clk), .Q(pipeline_PC_DX[30]), 
        .QN(n745) );
  DFF_X2 pipeline_PC_DX_reg_8_ ( .D(n5923), .CK(clk), .Q(pipeline_PC_DX[8]), 
        .QN(n723) );
  DFF_X2 pipeline_PC_DX_reg_7_ ( .D(n5925), .CK(clk), .Q(pipeline_PC_DX[7]), 
        .QN(n722) );
  DFF_X2 pipeline_PC_DX_reg_6_ ( .D(n5927), .CK(clk), .Q(pipeline_PC_DX[6]), 
        .QN(n721) );
  DFF_X2 pipeline_PC_DX_reg_5_ ( .D(n5929), .CK(clk), .Q(pipeline_PC_DX[5]), 
        .QN(n720) );
  DFF_X2 pipeline_PC_DX_reg_1_ ( .D(n5937), .CK(clk), .Q(pipeline_PC_DX[1]), 
        .QN(n716) );
  DFF_X2 pipeline_PC_DX_reg_0_ ( .D(n5939), .CK(clk), .Q(pipeline_PC_DX[0]), 
        .QN(n715) );
  DFF_X2 pipeline_PC_DX_reg_31_ ( .D(n5877), .CK(clk), .Q(pipeline_PC_DX[31]), 
        .QN(n746) );
  DFF_X2 pipeline_PC_IF_reg_10_ ( .D(n5961), .CK(clk), .QN(n12500) );
  DFF_X2 pipeline_csr_mepc_reg_1_ ( .D(n5874), .CK(clk), .QN(n1484) );
  DFF_X2 pipeline_csr_mepc_reg_0_ ( .D(n5875), .CK(clk), .QN(n1483) );
  DFF_X2 pipeline_csr_rdata_WB_reg_31_ ( .D(n6365), .CK(clk), .QN(n470) );
  DFF_X2 pipeline_csr_rdata_WB_reg_18_ ( .D(n6352), .CK(clk), .QN(n444) );
  DFF_X2 pipeline_csr_rdata_WB_reg_3_ ( .D(n6337), .CK(clk), .QN(n414) );
  DFF_X2 pipeline_csr_rdata_WB_reg_5_ ( .D(n6339), .CK(clk), .QN(n418) );
  DFF_X2 pipeline_PC_WB_reg_1_ ( .D(n5936), .CK(clk), .Q(n12383), .QN(n536) );
  DFF_X2 pipeline_PC_WB_reg_0_ ( .D(n5938), .CK(clk), .Q(n12616), .QN(n535) );
  DFF_X2 pipeline_csr_rdata_WB_reg_7_ ( .D(n6341), .CK(clk), .QN(n422) );
  DFF_X2 pipeline_csr_rdata_WB_reg_30_ ( .D(n6364), .CK(clk), .QN(n468) );
  DFF_X2 pipeline_csr_rdata_WB_reg_29_ ( .D(n6363), .CK(clk), .QN(n466) );
  DFF_X2 pipeline_csr_rdata_WB_reg_22_ ( .D(n6356), .CK(clk), .QN(n452) );
  DFF_X2 pipeline_csr_rdata_WB_reg_21_ ( .D(n6355), .CK(clk), .QN(n450) );
  DFF_X2 pipeline_csr_rdata_WB_reg_19_ ( .D(n6353), .CK(clk), .QN(n446) );
  DFF_X2 pipeline_csr_rdata_WB_reg_17_ ( .D(n6351), .CK(clk), .QN(n442) );
  DFF_X2 pipeline_csr_rdata_WB_reg_16_ ( .D(n6350), .CK(clk), .QN(n440) );
  DFF_X2 pipeline_csr_rdata_WB_reg_14_ ( .D(n6348), .CK(clk), .QN(n436) );
  DFF_X2 pipeline_csr_rdata_WB_reg_13_ ( .D(n6347), .CK(clk), .QN(n434) );
  DFF_X2 pipeline_csr_rdata_WB_reg_12_ ( .D(n6346), .CK(clk), .QN(n432) );
  DFF_X2 pipeline_csr_rdata_WB_reg_11_ ( .D(n6345), .CK(clk), .QN(n430) );
  DFF_X2 pipeline_csr_rdata_WB_reg_10_ ( .D(n6344), .CK(clk), .QN(n428) );
  DFF_X2 pipeline_csr_rdata_WB_reg_9_ ( .D(n6343), .CK(clk), .QN(n426) );
  DFF_X2 pipeline_csr_rdata_WB_reg_6_ ( .D(n6340), .CK(clk), .QN(n420) );
  DFF_X2 pipeline_csr_rdata_WB_reg_2_ ( .D(n6336), .CK(clk), .QN(n412) );
  DFF_X2 pipeline_csr_rdata_WB_reg_4_ ( .D(n6338), .CK(clk), .QN(n416) );
  DFF_X2 pipeline_csr_rdata_WB_reg_1_ ( .D(n6335), .CK(clk), .QN(n410) );
  DFF_X2 pipeline_csr_rdata_WB_reg_0_ ( .D(n6334), .CK(clk), .QN(n408) );
  DFF_X2 pipeline_csr_rdata_WB_reg_8_ ( .D(n6342), .CK(clk), .QN(n424) );
  DFF_X2 pipeline_csr_rdata_WB_reg_28_ ( .D(n6362), .CK(clk), .QN(n464) );
  DFF_X2 pipeline_csr_rdata_WB_reg_20_ ( .D(n6354), .CK(clk), .QN(n448) );
  DFF_X2 pipeline_csr_rdata_WB_reg_15_ ( .D(n6349), .CK(clk), .QN(n438) );
  DFF_X2 pipeline_csr_rdata_WB_reg_27_ ( .D(n6361), .CK(clk), .QN(n462) );
  DFF_X2 pipeline_csr_rdata_WB_reg_26_ ( .D(n6360), .CK(clk), .QN(n460) );
  DFF_X2 pipeline_csr_rdata_WB_reg_25_ ( .D(n6359), .CK(clk), .QN(n458) );
  DFF_X2 pipeline_csr_rdata_WB_reg_24_ ( .D(n6358), .CK(clk), .QN(n456) );
  DFF_X2 pipeline_csr_rdata_WB_reg_23_ ( .D(n6357), .CK(clk), .QN(n454) );
  DFF_X2 pipeline_store_data_WB_reg_11_ ( .D(n6321), .CK(clk), .Q(n13073), 
        .QN(n514) );
  DFF_X2 pipeline_store_data_WB_reg_8_ ( .D(n6324), .CK(clk), .Q(n13086), .QN(
        n511) );
  DFF_X2 pipeline_store_data_WB_reg_10_ ( .D(n6322), .CK(clk), .Q(n13072), 
        .QN(n513) );
  DFF_X2 pipeline_store_data_WB_reg_9_ ( .D(n6323), .CK(clk), .Q(n13088), .QN(
        n512) );
  DFF_X2 pipeline_store_data_WB_reg_16_ ( .D(n6316), .CK(clk), .Q(n13078), 
        .QN(n519) );
  DFF_X2 pipeline_store_data_WB_reg_19_ ( .D(n6313), .CK(clk), .Q(n13081), 
        .QN(n522) );
  DFF_X2 pipeline_store_data_WB_reg_18_ ( .D(n6314), .CK(clk), .Q(n13080), 
        .QN(n521) );
  DFF_X2 pipeline_store_data_WB_reg_28_ ( .D(n6304), .CK(clk), .Q(n13092), 
        .QN(n531) );
  DFF_X2 pipeline_store_data_WB_reg_13_ ( .D(n6319), .CK(clk), .Q(n13075), 
        .QN(n516) );
  DFF_X2 pipeline_store_data_WB_reg_14_ ( .D(n6318), .CK(clk), .Q(n13076), 
        .QN(n517) );
  DFF_X2 pipeline_store_data_WB_reg_23_ ( .D(n6309), .CK(clk), .Q(n13085), 
        .QN(n526) );
  DFF_X2 pipeline_store_data_WB_reg_29_ ( .D(n6303), .CK(clk), .Q(n13093), 
        .QN(n532) );
  DFF_X2 pipeline_store_data_WB_reg_30_ ( .D(n6302), .CK(clk), .Q(n13094), 
        .QN(n533) );
  DFF_X2 pipeline_store_data_WB_reg_12_ ( .D(n6320), .CK(clk), .Q(n13074), 
        .QN(n515) );
  DFF_X2 pipeline_store_data_WB_reg_15_ ( .D(n6317), .CK(clk), .Q(n13077), 
        .QN(n518) );
  DFF_X2 pipeline_store_data_WB_reg_27_ ( .D(n6305), .CK(clk), .Q(n13091), 
        .QN(n530) );
  DFF_X2 pipeline_store_data_WB_reg_25_ ( .D(n6307), .CK(clk), .Q(n13089), 
        .QN(n528) );
  DFF_X2 pipeline_store_data_WB_reg_22_ ( .D(n6310), .CK(clk), .Q(n13084), 
        .QN(n525) );
  DFF_X2 pipeline_store_data_WB_reg_21_ ( .D(n6311), .CK(clk), .Q(n13083), 
        .QN(n524) );
  DFF_X2 pipeline_store_data_WB_reg_26_ ( .D(n6306), .CK(clk), .Q(n13090), 
        .QN(n529) );
  DFF_X2 pipeline_store_data_WB_reg_17_ ( .D(n6315), .CK(clk), .Q(n13079), 
        .QN(n520) );
  DFF_X2 pipeline_store_data_WB_reg_24_ ( .D(n6308), .CK(clk), .Q(n13087), 
        .QN(n527) );
  DFF_X2 pipeline_store_data_WB_reg_20_ ( .D(n6312), .CK(clk), .Q(n13082), 
        .QN(n523) );
  DFF_X2 pipeline_ctrl_prev_killed_WB_reg ( .D(n6048), .CK(clk), .QN(n793) );
  DFF_X2 pipeline_ctrl_uses_md_WB_reg ( .D(n6251), .CK(clk), .Q(n9607), .QN(
        n787) );
  DFF_X2 pipeline_ctrl_store_in_WB_reg ( .D(n6253), .CK(clk), .Q(n9673), .QN(
        n790) );
  DFF_X2 pipeline_md_op_reg_1_ ( .D(n6242), .CK(clk), .Q(n10150), .QN(n964) );
  DFF_X2 pipeline_csr_mepc_reg_4_ ( .D(n5871), .CK(clk), .QN(n1487) );
  DFF_X2 pipeline_csr_mepc_reg_3_ ( .D(n5872), .CK(clk), .Q(n10496), .QN(n1486) );
  DFF_X2 pipeline_csr_mecode_reg_3_ ( .D(n5972), .CK(clk), .QN(n1482) );
  DFF_X2 pipeline_csr_to_host_reg_4_ ( .D(n6085), .CK(clk), .Q(n11237), .QN(
        n1259) );
  DFF_X2 pipeline_csr_mscratch_reg_4_ ( .D(n6140), .CK(clk), .Q(n11239), .QN(
        n1165) );
  DFF_X2 pipeline_csr_mie_reg_4_ ( .D(n6211), .CK(clk), .QN(n1519) );
  DFF_X2 pipeline_csr_mie_reg_30_ ( .D(n6237), .CK(clk), .Q(n9576), .QN(n1545)
         );
  DFF_X2 pipeline_csr_mie_reg_29_ ( .D(n6236), .CK(clk), .Q(n9575), .QN(n1544)
         );
  DFF_X2 pipeline_csr_mie_reg_27_ ( .D(n6234), .CK(clk), .Q(n9548), .QN(n1542)
         );
  DFF_X2 pipeline_csr_mie_reg_26_ ( .D(n6233), .CK(clk), .Q(n9554), .QN(n1541)
         );
  DFF_X2 pipeline_csr_mie_reg_25_ ( .D(n6232), .CK(clk), .Q(n9552), .QN(n1540)
         );
  DFF_X2 pipeline_csr_mie_reg_24_ ( .D(n6231), .CK(clk), .Q(n9553), .QN(n1539)
         );
  DFF_X2 pipeline_csr_mie_reg_23_ ( .D(n6230), .CK(clk), .Q(n9537), .QN(n1538)
         );
  DFF_X2 pipeline_csr_mie_reg_22_ ( .D(n6229), .CK(clk), .Q(n9571), .QN(n1537)
         );
  DFF_X2 pipeline_csr_mie_reg_21_ ( .D(n6228), .CK(clk), .Q(n9570), .QN(n1536)
         );
  DFF_X2 pipeline_csr_mie_reg_20_ ( .D(n6227), .CK(clk), .Q(n10896), .QN(n1535) );
  DFF_X2 pipeline_csr_mie_reg_19_ ( .D(n6226), .CK(clk), .Q(n9562), .QN(n1534)
         );
  DFF_X2 pipeline_csr_mie_reg_17_ ( .D(n6224), .CK(clk), .Q(n9563), .QN(n1532)
         );
  DFF_X2 pipeline_csr_mie_reg_16_ ( .D(n6223), .CK(clk), .Q(n9564), .QN(n1531)
         );
  DFF_X2 pipeline_csr_mie_reg_15_ ( .D(n6222), .CK(clk), .Q(n11114), .QN(n1530) );
  DFF_X2 pipeline_csr_mie_reg_14_ ( .D(n6221), .CK(clk), .Q(n9565), .QN(n1529)
         );
  DFF_X2 pipeline_csr_mie_reg_9_ ( .D(n6216), .CK(clk), .Q(n9536), .QN(n1524)
         );
  DFF_X2 pipeline_csr_mie_reg_6_ ( .D(n6213), .CK(clk), .Q(n10727), .QN(n1521)
         );
  DFF_X2 pipeline_csr_mie_reg_28_ ( .D(n6235), .CK(clk), .Q(n9577), .QN(n1543)
         );
  DFF_X2 pipeline_csr_mscratch_reg_3_ ( .D(n6141), .CK(clk), .QN(n1164) );
  DFF_X2 pipeline_csr_mie_reg_3_ ( .D(n6210), .CK(clk), .Q(n9547), .QN(n1518)
         );
  DFF_X2 pipeline_csr_mie_reg_5_ ( .D(n6212), .CK(clk), .QN(n1520) );
  DFF_X2 pipeline_csr_to_host_reg_30_ ( .D(n6111), .CK(clk), .Q(n10245), .QN(
        n1285) );
  DFF_X2 pipeline_csr_to_host_reg_29_ ( .D(n6110), .CK(clk), .Q(n10364), .QN(
        n1284) );
  DFF_X2 pipeline_csr_to_host_reg_27_ ( .D(n6108), .CK(clk), .Q(n10467), .QN(
        n1282) );
  DFF_X2 pipeline_csr_to_host_reg_26_ ( .D(n6107), .CK(clk), .Q(n10543), .QN(
        n1281) );
  DFF_X2 pipeline_csr_to_host_reg_25_ ( .D(n6106), .CK(clk), .Q(n10597), .QN(
        n1280) );
  DFF_X2 pipeline_csr_to_host_reg_24_ ( .D(n6105), .CK(clk), .Q(n10651), .QN(
        n1279) );
  DFF_X2 pipeline_csr_to_host_reg_23_ ( .D(n6104), .CK(clk), .Q(n10705), .QN(
        n1278) );
  DFF_X2 pipeline_csr_to_host_reg_22_ ( .D(n6103), .CK(clk), .Q(n10756), .QN(
        n1277) );
  DFF_X2 pipeline_csr_to_host_reg_21_ ( .D(n6102), .CK(clk), .Q(n10841), .QN(
        n1276) );
  DFF_X2 pipeline_csr_to_host_reg_20_ ( .D(n6101), .CK(clk), .QN(n1275) );
  DFF_X2 pipeline_csr_to_host_reg_19_ ( .D(n6100), .CK(clk), .Q(n10949), .QN(
        n1274) );
  DFF_X2 pipeline_csr_to_host_reg_18_ ( .D(n6099), .CK(clk), .QN(n1273) );
  DFF_X2 pipeline_csr_to_host_reg_17_ ( .D(n6098), .CK(clk), .Q(n11056), .QN(
        n1272) );
  DFF_X2 pipeline_csr_to_host_reg_16_ ( .D(n6097), .CK(clk), .Q(n11083), .QN(
        n1271) );
  DFF_X2 pipeline_csr_to_host_reg_15_ ( .D(n6096), .CK(clk), .QN(n1270) );
  DFF_X2 pipeline_csr_to_host_reg_14_ ( .D(n6095), .CK(clk), .Q(n11141), .QN(
        n1269) );
  DFF_X2 pipeline_csr_to_host_reg_13_ ( .D(n6094), .CK(clk), .Q(n11029), .QN(
        n1268) );
  DFF_X2 pipeline_csr_to_host_reg_12_ ( .D(n6093), .CK(clk), .Q(n10868), .QN(
        n1267) );
  DFF_X2 pipeline_csr_to_host_reg_11_ ( .D(n6092), .CK(clk), .Q(n10922), .QN(
        n1266) );
  DFF_X2 pipeline_csr_to_host_reg_10_ ( .D(n6091), .CK(clk), .Q(n10976), .QN(
        n1265) );
  DFF_X2 pipeline_csr_to_host_reg_9_ ( .D(n6090), .CK(clk), .Q(n10570), .QN(
        n1264) );
  DFF_X2 pipeline_csr_to_host_reg_6_ ( .D(n6087), .CK(clk), .Q(n10730), .QN(
        n1261) );
  DFF_X2 pipeline_csr_from_host_reg_20_ ( .D(n6061), .CK(clk), .QN(n1243) );
  DFF_X2 pipeline_csr_from_host_reg_15_ ( .D(n6066), .CK(clk), .QN(n1238) );
  DFF_X2 pipeline_csr_from_host_reg_6_ ( .D(n6075), .CK(clk), .Q(n10729), .QN(
        n1229) );
  DFF_X2 pipeline_csr_to_host_reg_28_ ( .D(n6109), .CK(clk), .QN(n1283) );
  DFF_X2 pipeline_csr_to_host_reg_5_ ( .D(n6086), .CK(clk), .Q(n10780), .QN(
        n1260) );
  DFF_X2 pipeline_csr_mscratch_reg_5_ ( .D(n6139), .CK(clk), .QN(n1166) );
  DFF_X2 pipeline_csr_to_host_reg_31_ ( .D(n6367), .CK(clk), .Q(n10289), .QN(
        n1286) );
  DFF_X2 pipeline_csr_mint_reg ( .D(n5983), .CK(clk), .Q(n10286), .QN(n1478)
         );
  DFF_X2 pipeline_csr_mepc_reg_2_ ( .D(n5873), .CK(clk), .Q(n10406), .QN(n1485) );
  DFF_X2 pipeline_csr_mecode_reg_2_ ( .D(n5973), .CK(clk), .QN(n1481) );
  DFF_X2 pipeline_csr_mepc_reg_26_ ( .D(n5849), .CK(clk), .Q(n10540), .QN(
        n1509) );
  DFF_X2 pipeline_csr_mepc_reg_25_ ( .D(n5850), .CK(clk), .Q(n10594), .QN(
        n1508) );
  DFF_X2 pipeline_csr_mepc_reg_24_ ( .D(n5851), .CK(clk), .Q(n10648), .QN(
        n1507) );
  DFF_X2 pipeline_csr_mepc_reg_23_ ( .D(n5852), .CK(clk), .Q(n10702), .QN(
        n1506) );
  DFF_X2 pipeline_csr_mepc_reg_22_ ( .D(n5853), .CK(clk), .Q(n10753), .QN(
        n1505) );
  DFF_X2 pipeline_csr_mepc_reg_21_ ( .D(n5854), .CK(clk), .Q(n10838), .QN(
        n1504) );
  DFF_X2 pipeline_csr_mepc_reg_20_ ( .D(n5855), .CK(clk), .QN(n1503) );
  DFF_X2 pipeline_csr_mepc_reg_19_ ( .D(n5856), .CK(clk), .Q(n10946), .QN(
        n1502) );
  DFF_X2 pipeline_csr_mepc_reg_18_ ( .D(n5857), .CK(clk), .QN(n1501) );
  DFF_X2 pipeline_csr_mepc_reg_17_ ( .D(n5858), .CK(clk), .Q(n11053), .QN(
        n1500) );
  DFF_X2 pipeline_csr_mepc_reg_16_ ( .D(n5859), .CK(clk), .Q(n11080), .QN(
        n1499) );
  DFF_X2 pipeline_csr_mepc_reg_15_ ( .D(n5860), .CK(clk), .QN(n1498) );
  DFF_X2 pipeline_csr_mepc_reg_14_ ( .D(n5861), .CK(clk), .Q(n11137), .QN(
        n1497) );
  DFF_X2 pipeline_csr_mepc_reg_13_ ( .D(n5862), .CK(clk), .Q(n11026), .QN(
        n1496) );
  DFF_X2 pipeline_csr_mepc_reg_12_ ( .D(n5863), .CK(clk), .Q(n10865), .QN(
        n1495) );
  DFF_X2 pipeline_csr_mepc_reg_11_ ( .D(n5864), .CK(clk), .Q(n10919), .QN(
        n1494) );
  DFF_X2 pipeline_csr_mepc_reg_10_ ( .D(n5865), .CK(clk), .Q(n10973), .QN(
        n1493) );
  DFF_X2 pipeline_csr_mepc_reg_9_ ( .D(n5866), .CK(clk), .Q(n10567), .QN(n1492) );
  DFF_X2 pipeline_csr_mepc_reg_6_ ( .D(n5869), .CK(clk), .QN(n1489) );
  DFF_X2 pipeline_csr_mepc_reg_5_ ( .D(n5870), .CK(clk), .Q(n10781), .QN(n1488) );
  DFF_X2 pipeline_csr_to_host_reg_8_ ( .D(n6089), .CK(clk), .QN(n1263) );
  DFF_X2 pipeline_csr_from_host_reg_8_ ( .D(n6073), .CK(clk), .QN(n1231) );
  DFF_X2 pipeline_csr_to_host_reg_7_ ( .D(n6088), .CK(clk), .Q(n10679), .QN(
        n1262) );
  DFF_X2 pipeline_csr_mepc_reg_7_ ( .D(n5868), .CK(clk), .Q(n10676), .QN(n1490) );
  DFF_X2 pipeline_csr_to_host_reg_2_ ( .D(n6083), .CK(clk), .Q(n10403), .QN(
        n1257) );
  DFF_X2 pipeline_csr_mscratch_reg_2_ ( .D(n6142), .CK(clk), .QN(n1163) );
  DFF_X2 pipeline_csr_mie_reg_2_ ( .D(n6209), .CK(clk), .QN(n1517) );
  DFF_X2 pipeline_csr_to_host_reg_0_ ( .D(n6112), .CK(clk), .QN(n1255) );
  DFF_X2 pipeline_csr_mscratch_reg_0_ ( .D(n6144), .CK(clk), .Q(n11267), .QN(
        n1161) );
  DFF_X2 pipeline_csr_mie_reg_0_ ( .D(n6239), .CK(clk), .Q(n11271), .QN(n1515)
         );
  DFF_X2 pipeline_csr_mepc_reg_27_ ( .D(n5848), .CK(clk), .Q(n10464), .QN(
        n1510) );
  DFF_X2 pipeline_csr_mepc_reg_8_ ( .D(n5867), .CK(clk), .QN(n1491) );
  DFF_X2 pipeline_csr_mecode_reg_0_ ( .D(n5975), .CK(clk), .Q(n12627) );
  DFF_X2 pipeline_csr_mepc_reg_28_ ( .D(n5847), .CK(clk), .Q(n10429), .QN(
        n1511) );
  DFF_X2 pipeline_csr_mie_reg_1_ ( .D(n6208), .CK(clk), .QN(n1516) );
  DFF_X2 pipeline_csr_mepc_reg_29_ ( .D(n5846), .CK(clk), .Q(n10361), .QN(
        n1512) );
  DFF_X2 pipeline_csr_to_host_reg_1_ ( .D(n6082), .CK(clk), .QN(n1256) );
  DFF_X2 pipeline_csr_mscratch_reg_1_ ( .D(n6143), .CK(clk), .Q(n10322), .QN(
        n1162) );
  DFF_X2 pipeline_csr_mepc_reg_30_ ( .D(n5845), .CK(clk), .Q(n10241), .QN(
        n1513) );
  DFF_X2 pipeline_csr_mepc_reg_31_ ( .D(n5844), .CK(clk), .Q(n10285), .QN(
        n1514) );
  DFF_X2 pipeline_csr_mecode_reg_1_ ( .D(n5974), .CK(clk), .Q(n10321), .QN(
        n1480) );
  DFF_X2 pipeline_inst_DX_reg_8_ ( .D(n6265), .CK(clk), .Q(n10137), .QN(n595)
         );
  DFF_X2 pipeline_inst_DX_reg_7_ ( .D(n6263), .CK(clk), .Q(n10138), .QN(n594)
         );
  DFF_X2 pipeline_PC_IF_reg_25_ ( .D(n5946), .CK(clk), .QN(n12441) );
  DFF_X2 pipeline_PC_IF_reg_9_ ( .D(n5962), .CK(clk), .QN(n12504) );
  DFF_X2 pipeline_PC_IF_reg_29_ ( .D(n5942), .CK(clk), .QN(n12425) );
  DFF_X2 pipeline_PC_IF_reg_28_ ( .D(n5943), .CK(clk), .QN(n12429) );
  DFF_X2 pipeline_PC_IF_reg_26_ ( .D(n5945), .CK(clk), .QN(n12437) );
  DFF_X2 pipeline_PC_IF_reg_24_ ( .D(n5947), .CK(clk), .QN(n12445) );
  DFF_X2 pipeline_PC_IF_reg_23_ ( .D(n5948), .CK(clk), .QN(n12449) );
  DFF_X2 pipeline_PC_IF_reg_31_ ( .D(n5940), .CK(clk), .QN(n12416) );
  DFF_X2 pipeline_PC_IF_reg_30_ ( .D(n5941), .CK(clk), .QN(n12421) );
  DFF_X2 pipeline_PC_IF_reg_19_ ( .D(n5952), .CK(clk), .QN(n12465) );
  DFF_X2 pipeline_PC_IF_reg_27_ ( .D(n5944), .CK(clk), .QN(n12433) );
  DFF_X2 pipeline_PC_IF_reg_22_ ( .D(n5949), .CK(clk), .QN(n12453) );
  DFF_X2 pipeline_PC_IF_reg_18_ ( .D(n5953), .CK(clk), .QN(n12469) );
  DFF_X2 pipeline_PC_IF_reg_21_ ( .D(n5950), .CK(clk), .QN(n12457) );
  DFF_X2 pipeline_PC_IF_reg_20_ ( .D(n5951), .CK(clk), .QN(n12461) );
  NOR2_X2 U6281 ( .A1(n12493), .A2(n9485), .ZN(n12494) );
  BUF_X2 U6282 ( .A(pipeline_alu_src_a[13]), .Z(n6566) );
  NOR2_X2 U6283 ( .A1(n12599), .A2(n6944), .ZN(n9613) );
  OAI221_X2 U6284 ( .B1(n9802), .B2(n9448), .C1(n9632), .C2(n9396), .A(n10043), 
        .ZN(n6556) );
  OAI221_X2 U6285 ( .B1(n9802), .B2(n9448), .C1(n9632), .C2(n9396), .A(n10043), 
        .ZN(n6557) );
  INV_X8 U6286 ( .A(n8232), .ZN(n8257) );
  NAND2_X4 U6287 ( .A1(n7192), .A2(n7163), .ZN(n11318) );
  NAND2_X4 U6288 ( .A1(n7192), .A2(n9402), .ZN(n12612) );
  NAND2_X4 U6289 ( .A1(n11323), .A2(n13130), .ZN(n3683) );
  NAND4_X4 U6290 ( .A1(n10334), .A2(n10336), .A3(n9402), .A4(n6711), .ZN(
        n12255) );
  NAND2_X4 U6291 ( .A1(n7190), .A2(n10351), .ZN(n12352) );
  NAND2_X4 U6292 ( .A1(n10520), .A2(n10519), .ZN(n12347) );
  NAND2_X4 U6293 ( .A1(n7190), .A2(n10518), .ZN(n12349) );
  AOI21_X4 U6294 ( .B1(n9468), .B2(n10343), .A(n11198), .ZN(n9403) );
  NAND2_X4 U6295 ( .A1(n7016), .A2(n7075), .ZN(n11282) );
  INV_X8 U6296 ( .A(n8250), .ZN(n8253) );
  INV_X4 U6297 ( .A(n8250), .ZN(n8252) );
  OAI221_X2 U6298 ( .B1(n597), .B2(n9795), .C1(n9707), .C2(n10056), .A(n9706), 
        .ZN(n9339) );
  INV_X8 U6299 ( .A(n9303), .ZN(n9328) );
  AND4_X2 U6300 ( .A1(n8143), .A2(n8144), .A3(n8145), .A4(n8146), .ZN(n7135)
         );
  OAI221_X4 U6301 ( .B1(n9487), .B2(n12516), .C1(n1489), .C2(n6661), .A(n12515), .ZN(pipeline_PCmux_base[6]) );
  OAI21_X4 U6302 ( .B1(n10014), .B2(n10013), .A(n10012), .ZN(n10024) );
  AOI21_X4 U6303 ( .B1(n9995), .B2(n9996), .A(n9994), .ZN(n10014) );
  OAI221_X1 U6304 ( .B1(n9488), .B2(n12429), .C1(n1511), .C2(n6661), .A(n12428), .ZN(pipeline_PCmux_base[28]) );
  INV_X4 U6305 ( .A(pipeline_alu_src_a[26]), .ZN(n6558) );
  INV_X4 U6306 ( .A(n6558), .ZN(n6559) );
  INV_X4 U6307 ( .A(n6558), .ZN(n6560) );
  INV_X4 U6308 ( .A(n6558), .ZN(n6561) );
  AND4_X2 U6309 ( .A1(n7313), .A2(n7314), .A3(n7315), .A4(n7316), .ZN(n7148)
         );
  NAND2_X4 U6310 ( .A1(n9391), .A2(n10258), .ZN(n9338) );
  AOI221_X2 U6311 ( .B1(pipeline_PC_DX[11]), .B2(n9337), .C1(
        pipeline_handler_PC[11]), .C2(n6630), .A(n12494), .ZN(n12495) );
  INV_X1 U6312 ( .A(n12599), .ZN(n12149) );
  AOI21_X4 U6313 ( .B1(n10054), .B2(n10053), .A(n10052), .ZN(n10069) );
  OAI21_X4 U6314 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10053) );
  INV_X4 U6315 ( .A(pipeline_alu_src_a[28]), .ZN(n6562) );
  INV_X4 U6316 ( .A(n6562), .ZN(n6563) );
  INV_X4 U6317 ( .A(n6562), .ZN(n6564) );
  INV_X4 U6318 ( .A(n6562), .ZN(n6565) );
  NOR2_X1 U6319 ( .A1(n12426), .A2(n9484), .ZN(n12427) );
  NAND2_X4 U6320 ( .A1(n12561), .A2(n12557), .ZN(n9337) );
  BUF_X4 U6321 ( .A(pipeline_alu_src_a[13]), .Z(n6567) );
  BUF_X4 U6322 ( .A(pipeline_alu_src_a[13]), .Z(n6568) );
  NAND2_X1 U6323 ( .A1(n9914), .A2(n9860), .ZN(n9919) );
  INV_X4 U6324 ( .A(pipeline_alu_src_a[10]), .ZN(n6569) );
  INV_X4 U6325 ( .A(n6569), .ZN(n6570) );
  INV_X1 U6326 ( .A(n6569), .ZN(n6571) );
  INV_X1 U6327 ( .A(n6569), .ZN(n6572) );
  INV_X4 U6328 ( .A(pipeline_rs2_data_bypassed[4]), .ZN(n9792) );
  OAI22_X2 U6329 ( .A1(n9847), .A2(n9448), .B1(n10236), .B2(n9915), .ZN(
        pipeline_alu_src_b[7]) );
  OAI221_X2 U6330 ( .B1(n9931), .B2(n10056), .C1(n602), .C2(n9397), .A(n9967), 
        .ZN(pipeline_alu_src_b[13]) );
  OAI221_X2 U6331 ( .B1(n9833), .B2(n10056), .C1(n603), .C2(n10044), .A(n9967), 
        .ZN(pipeline_alu_src_b[14]) );
  OAI221_X2 U6332 ( .B1(n10045), .B2(n9448), .C1(n713), .C2(n10044), .A(n10043), .ZN(pipeline_alu_src_b[30]) );
  AOI221_X2 U6333 ( .B1(pipeline_PC_DX[15]), .B2(n9336), .C1(
        pipeline_handler_PC[15]), .C2(n6630), .A(n12478), .ZN(n12479) );
  NOR2_X2 U6334 ( .A1(n12477), .A2(n9485), .ZN(n12478) );
  OAI221_X2 U6335 ( .B1(n9488), .B2(n12473), .C1(n1500), .C2(n6661), .A(n12472), .ZN(pipeline_PCmux_base[17]) );
  NAND3_X2 U6336 ( .A1(n6967), .A2(n6968), .A3(n12475), .ZN(
        pipeline_PCmux_base[16]) );
  INV_X4 U6337 ( .A(n9338), .ZN(n6942) );
  INV_X4 U6338 ( .A(pipeline_alu_src_b[7]), .ZN(n11885) );
  OAI22_X2 U6339 ( .A1(n730), .A2(n9445), .B1(n12477), .B2(n9443), .ZN(
        pipeline_alu_src_a[15]) );
  OAI22_X2 U6340 ( .A1(n743), .A2(n9445), .B1(n12426), .B2(n9443), .ZN(
        pipeline_alu_src_a[28]) );
  NAND2_X2 U6341 ( .A1(n6742), .A2(n12403), .ZN(n12411) );
  INV_X4 U6342 ( .A(pipeline_regfile_N18), .ZN(n9658) );
  NAND2_X2 U6343 ( .A1(n9389), .A2(n9390), .ZN(n9391) );
  AOI21_X2 U6344 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(n10348) );
  NAND2_X2 U6345 ( .A1(n9724), .A2(n9723), .ZN(n9393) );
  OAI22_X2 U6346 ( .A1(n725), .A2(n9445), .B1(n12497), .B2(n9443), .ZN(
        pipeline_alu_src_a[10]) );
  OAI221_X2 U6347 ( .B1(n9802), .B2(n9448), .C1(n9632), .C2(n9396), .A(n10043), 
        .ZN(pipeline_alu_src_b[29]) );
  OAI22_X2 U6348 ( .A1(n7061), .A2(n7139), .B1(n12941), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[8]) );
  OAI22_X2 U6349 ( .A1(n7061), .A2(n7100), .B1(n12904), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[15]) );
  NAND3_X2 U6350 ( .A1(n7058), .A2(n7059), .A3(n7060), .ZN(dmem_haddr[31]) );
  NAND3_X2 U6351 ( .A1(n9801), .A2(n10081), .A3(n6578), .ZN(n6573) );
  AND2_X4 U6352 ( .A1(n12660), .A2(n12659), .ZN(n6574) );
  AND3_X4 U6353 ( .A1(n12994), .A2(n9668), .A3(n9669), .ZN(n6575) );
  AND2_X4 U6354 ( .A1(n7259), .A2(n7260), .ZN(n6576) );
  OR2_X2 U6355 ( .A1(n12474), .A2(n9485), .ZN(n6577) );
  NAND2_X2 U6356 ( .A1(n11404), .A2(n11405), .ZN(n12565) );
  AND2_X4 U6357 ( .A1(n10074), .A2(n9693), .ZN(n6578) );
  INV_X4 U6358 ( .A(n7050), .ZN(n8271) );
  NAND3_X2 U6359 ( .A1(pipeline_regfile_N19), .A2(n693), .A3(n9658), .ZN(n7050) );
  NAND2_X2 U6360 ( .A1(n637), .A2(n6579), .ZN(n6710) );
  NOR2_X2 U6361 ( .A1(n636), .A2(n638), .ZN(n6579) );
  INV_X8 U6362 ( .A(n6710), .ZN(n9321) );
  NAND2_X2 U6363 ( .A1(n7003), .A2(n693), .ZN(n6580) );
  INV_X4 U6364 ( .A(n12542), .ZN(n9481) );
  AOI221_X1 U6365 ( .B1(pipeline_md_N58), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[29]), .A(n10377), .ZN(n10378) );
  AOI221_X1 U6366 ( .B1(n9471), .B2(n12064), .C1(n12276), .C2(n9334), .A(
        n11169), .ZN(n11757) );
  OR2_X1 U6367 ( .A1(n8502), .A2(n8278), .ZN(n6581) );
  OR2_X1 U6368 ( .A1(n8503), .A2(n9306), .ZN(n6582) );
  NAND2_X2 U6369 ( .A1(n6581), .A2(n6582), .ZN(n8501) );
  AND2_X2 U6370 ( .A1(pipeline_PC_DX[4]), .A2(n6958), .ZN(n6583) );
  AND2_X1 U6371 ( .A1(pipeline_handler_PC[4]), .A2(n6630), .ZN(n6584) );
  NOR3_X1 U6372 ( .A1(n6583), .A2(n6584), .A3(n12523), .ZN(n12524) );
  NOR2_X1 U6373 ( .A1(n12522), .A2(n9486), .ZN(n12523) );
  OR2_X1 U6374 ( .A1(n9387), .A2(n9455), .ZN(n6585) );
  OR2_X1 U6375 ( .A1(n9334), .A2(n9451), .ZN(n6586) );
  NAND2_X2 U6376 ( .A1(n6585), .A2(n6586), .ZN(n9858) );
  NOR2_X1 U6377 ( .A1(n9856), .A2(n9858), .ZN(n9862) );
  AND2_X4 U6378 ( .A1(pipeline_PC_DX[20]), .A2(n9482), .ZN(n6587) );
  AND2_X1 U6379 ( .A1(pipeline_handler_PC[20]), .A2(n6630), .ZN(n6588) );
  NOR3_X1 U6380 ( .A1(n6587), .A2(n6588), .A3(n12459), .ZN(n12460) );
  NOR2_X1 U6381 ( .A1(n12458), .A2(n9484), .ZN(n12459) );
  NAND2_X2 U6382 ( .A1(n12662), .A2(n12661), .ZN(n6589) );
  NAND2_X2 U6383 ( .A1(pipeline_alu_N89), .A2(n6813), .ZN(n6590) );
  AND3_X2 U6384 ( .A1(n6589), .A2(n6590), .A3(n6574), .ZN(n12663) );
  NAND2_X2 U6385 ( .A1(n12664), .A2(n12663), .ZN(dmem_haddr[30]) );
  NAND2_X2 U6386 ( .A1(pipeline_regfile_data[353]), .A2(n8249), .ZN(n6591) );
  NAND2_X1 U6387 ( .A1(pipeline_regfile_data[289]), .A2(n8253), .ZN(n6592) );
  AND3_X2 U6388 ( .A1(n6591), .A2(n6592), .A3(n6576), .ZN(n7258) );
  OR2_X1 U6389 ( .A1(n9487), .A2(n12534), .ZN(n6593) );
  OR2_X1 U6390 ( .A1(n1485), .A2(n6661), .ZN(n6594) );
  NAND3_X2 U6391 ( .A1(n6593), .A2(n6594), .A3(n12533), .ZN(
        pipeline_PCmux_base[2]) );
  AOI221_X1 U6392 ( .B1(pipeline_PC_DX[2]), .B2(n9480), .C1(
        pipeline_handler_PC[2]), .C2(n6630), .A(n12531), .ZN(n12533) );
  AND2_X2 U6393 ( .A1(n7352), .A2(n7353), .ZN(n7351) );
  OAI22_X2 U6394 ( .A1(n722), .A2(n9445), .B1(n12509), .B2(n9443), .ZN(
        pipeline_alu_src_a[7]) );
  AND2_X2 U6395 ( .A1(pipeline_regfile_data[836]), .A2(n6729), .ZN(n7376) );
  INV_X8 U6396 ( .A(n9370), .ZN(imem_haddr[24]) );
  NAND2_X1 U6397 ( .A1(n9386), .A2(n9389), .ZN(n9784) );
  OAI22_X1 U6398 ( .A1(n12449), .A2(n12632), .B1(n9372), .B2(n9493), .ZN(n5948) );
  INV_X8 U6399 ( .A(n9372), .ZN(imem_haddr[23]) );
  INV_X4 U6400 ( .A(pipeline_alu_src_a[15]), .ZN(n6595) );
  INV_X4 U6401 ( .A(n6595), .ZN(n6596) );
  INV_X1 U6402 ( .A(n6595), .ZN(n6597) );
  INV_X1 U6403 ( .A(n6595), .ZN(n6598) );
  INV_X4 U6404 ( .A(pipeline_alu_src_a[6]), .ZN(n6604) );
  OAI22_X2 U6405 ( .A1(n721), .A2(n9445), .B1(n12513), .B2(n9785), .ZN(
        pipeline_alu_src_a[6]) );
  INV_X4 U6406 ( .A(n9857), .ZN(n9856) );
  AND2_X2 U6407 ( .A1(n7264), .A2(n7265), .ZN(n7255) );
  AOI221_X2 U6408 ( .B1(pipeline_regfile_data[329]), .B2(n9324), .C1(
        pipeline_regfile_data[265]), .C2(n9327), .A(n8573), .ZN(n8568) );
  INV_X2 U6409 ( .A(n7375), .ZN(n7374) );
  AOI221_X1 U6410 ( .B1(pipeline_regfile_data[371]), .B2(n9309), .C1(
        pipeline_regfile_data[307]), .C2(n9316), .A(n8890), .ZN(n8889) );
  AOI221_X1 U6411 ( .B1(pipeline_regfile_data[112]), .B2(n9309), .C1(
        pipeline_regfile_data[48]), .C2(n9316), .A(n8802), .ZN(n8801) );
  AOI221_X1 U6412 ( .B1(pipeline_regfile_data[368]), .B2(n9309), .C1(
        pipeline_regfile_data[304]), .C2(n9316), .A(n8794), .ZN(n8793) );
  AOI221_X1 U6413 ( .B1(pipeline_regfile_data[109]), .B2(n9309), .C1(
        pipeline_regfile_data[45]), .C2(n9316), .A(n8706), .ZN(n8705) );
  AOI221_X1 U6414 ( .B1(pipeline_regfile_data[365]), .B2(n9309), .C1(
        pipeline_regfile_data[301]), .C2(n9316), .A(n8698), .ZN(n8697) );
  INV_X1 U6415 ( .A(n9481), .ZN(n9482) );
  INV_X4 U6416 ( .A(n9481), .ZN(n6969) );
  AND2_X2 U6417 ( .A1(n7480), .A2(n7481), .ZN(n7479) );
  NOR2_X1 U6418 ( .A1(pipeline_alu_src_b[26]), .A2(n12357), .ZN(n12088) );
  BUF_X4 U6419 ( .A(n8267), .Z(n6599) );
  INV_X1 U6420 ( .A(n6580), .ZN(n8267) );
  OAI221_X2 U6421 ( .B1(n598), .B2(n9795), .C1(n9792), .C2(n9448), .A(n9791), 
        .ZN(n6600) );
  OAI22_X1 U6422 ( .A1(n1483), .A2(n6661), .B1(n9488), .B2(n12539), .ZN(n12540) );
  AOI221_X1 U6423 ( .B1(pipeline_regfile_data[370]), .B2(n9309), .C1(
        pipeline_regfile_data[306]), .C2(n9313), .A(n8858), .ZN(n8857) );
  AOI221_X1 U6424 ( .B1(pipeline_regfile_data[369]), .B2(n9309), .C1(
        pipeline_regfile_data[305]), .C2(n9313), .A(n8826), .ZN(n8825) );
  INV_X2 U6425 ( .A(n9890), .ZN(n9873) );
  AND4_X2 U6426 ( .A1(n8753), .A2(n8754), .A3(n8755), .A4(n8756), .ZN(n7099)
         );
  INV_X4 U6427 ( .A(pipeline_alu_src_a[27]), .ZN(n6601) );
  INV_X1 U6428 ( .A(n6601), .ZN(n6602) );
  INV_X1 U6429 ( .A(n6601), .ZN(n6603) );
  INV_X1 U6430 ( .A(n6604), .ZN(n6605) );
  INV_X1 U6431 ( .A(n6604), .ZN(n6606) );
  INV_X4 U6432 ( .A(pipeline_alu_src_a[25]), .ZN(n6607) );
  INV_X4 U6433 ( .A(n6607), .ZN(n6608) );
  INV_X4 U6434 ( .A(n6607), .ZN(n6609) );
  INV_X4 U6435 ( .A(pipeline_alu_src_a[7]), .ZN(n6610) );
  INV_X1 U6436 ( .A(n6610), .ZN(n6611) );
  INV_X1 U6437 ( .A(n6610), .ZN(n6612) );
  INV_X4 U6438 ( .A(pipeline_alu_src_a[11]), .ZN(n6613) );
  INV_X1 U6439 ( .A(n6613), .ZN(n6614) );
  INV_X4 U6440 ( .A(pipeline_alu_src_b[0]), .ZN(n6615) );
  INV_X1 U6441 ( .A(n6615), .ZN(n6616) );
  INV_X4 U6442 ( .A(n6615), .ZN(n6617) );
  INV_X1 U6443 ( .A(n6615), .ZN(n6618) );
  OAI22_X2 U6444 ( .A1(n746), .A2(n9445), .B1(n12413), .B2(n9443), .ZN(
        pipeline_alu_N316) );
  AOI22_X2 U6445 ( .A1(n9981), .A2(n9980), .B1(n9979), .B2(n9978), .ZN(n9982)
         );
  INV_X4 U6446 ( .A(pipeline_alu_src_a[1]), .ZN(n6631) );
  OAI22_X2 U6447 ( .A1(n716), .A2(n9445), .B1(n6636), .B2(n9785), .ZN(
        pipeline_alu_src_a[1]) );
  OAI221_X2 U6448 ( .B1(n595), .B2(n9795), .C1(n9716), .C2(n9448), .A(n9715), 
        .ZN(pipeline_alu_src_b[1]) );
  OAI22_X2 U6449 ( .A1(n720), .A2(n9445), .B1(n12517), .B2(n9785), .ZN(
        pipeline_alu_src_a[5]) );
  INV_X4 U6450 ( .A(pipeline_rs1_data_bypassed[5]), .ZN(n12517) );
  OAI22_X2 U6451 ( .A1(n6633), .A2(n9454), .B1(n7009), .B2(n6744), .ZN(n9890)
         );
  NAND2_X2 U6452 ( .A1(n9311), .A2(n6736), .ZN(n9291) );
  AOI22_X2 U6453 ( .A1(n10011), .A2(n10010), .B1(n10009), .B2(n10008), .ZN(
        n10012) );
  OAI22_X2 U6454 ( .A1(n719), .A2(n9445), .B1(n12522), .B2(n9785), .ZN(n6928)
         );
  INV_X4 U6455 ( .A(pipeline_alu_src_a[2]), .ZN(n12274) );
  INV_X4 U6456 ( .A(n9483), .ZN(n9486) );
  OAI221_X2 U6457 ( .B1(n9488), .B2(n12469), .C1(n1501), .C2(n6661), .A(n12468), .ZN(pipeline_PCmux_base[18]) );
  OAI221_X2 U6458 ( .B1(n9488), .B2(n12453), .C1(n1505), .C2(n6661), .A(n12452), .ZN(pipeline_PCmux_base[22]) );
  OAI221_X2 U6459 ( .B1(n9488), .B2(n12465), .C1(n1502), .C2(n6661), .A(n12464), .ZN(pipeline_PCmux_base[19]) );
  NAND2_X2 U6460 ( .A1(n9561), .A2(n9560), .ZN(n9585) );
  NAND2_X2 U6461 ( .A1(n8446), .A2(n8447), .ZN(n8445) );
  BUF_X4 U6462 ( .A(n12994), .Z(n6941) );
  INV_X4 U6463 ( .A(n9291), .ZN(n8302) );
  OAI221_X2 U6464 ( .B1(n594), .B2(n9795), .C1(n9720), .C2(n10056), .A(n9719), 
        .ZN(pipeline_alu_src_b[0]) );
  AOI22_X2 U6465 ( .A1(pipeline_PC_DX[0]), .A2(n9446), .B1(
        pipeline_rs1_data_bypassed[0]), .B2(n9444), .ZN(n6943) );
  NAND2_X2 U6466 ( .A1(n6995), .A2(n6996), .ZN(pipeline_alu_src_a[17]) );
  INV_X4 U6467 ( .A(n6975), .ZN(n11405) );
  INV_X4 U6468 ( .A(n6943), .ZN(pipeline_alu_src_a[0]) );
  OAI221_X2 U6469 ( .B1(n9805), .B2(n9448), .C1(n8214), .C2(n9397), .A(n10043), 
        .ZN(pipeline_alu_src_b[24]) );
  OAI22_X2 U6470 ( .A1(n740), .A2(n9445), .B1(n12438), .B2(n9443), .ZN(
        pipeline_alu_src_a[25]) );
  OAI22_X2 U6471 ( .A1(n741), .A2(n9445), .B1(n12434), .B2(n9443), .ZN(
        pipeline_alu_src_a[26]) );
  INV_X4 U6472 ( .A(pipeline_rs1_data_bypassed[23]), .ZN(n12446) );
  AOI221_X1 U6473 ( .B1(pipeline_regfile_data[952]), .B2(n6728), .C1(
        pipeline_regfile_data[696]), .C2(n6720), .A(n7988), .ZN(n7987) );
  NAND2_X2 U6474 ( .A1(pipeline_regfile_data[689]), .A2(n6720), .ZN(n7000) );
  AOI22_X2 U6475 ( .A1(n6931), .A2(n9304), .B1(n6932), .B2(n6776), .ZN(n6930)
         );
  INV_X4 U6476 ( .A(n10783), .ZN(n13116) );
  NAND2_X2 U6477 ( .A1(n13144), .A2(n12846), .ZN(n4229) );
  OAI22_X2 U6478 ( .A1(n719), .A2(n9445), .B1(n12522), .B2(n9785), .ZN(n6927)
         );
  OAI22_X2 U6479 ( .A1(n726), .A2(n9445), .B1(n12493), .B2(n9443), .ZN(
        pipeline_alu_src_a[11]) );
  INV_X4 U6480 ( .A(pipeline_alu_src_a[17]), .ZN(n11546) );
  INV_X4 U6481 ( .A(n6780), .ZN(n9488) );
  INV_X4 U6482 ( .A(n13168), .ZN(n9372) );
  INV_X4 U6483 ( .A(n13167), .ZN(n9370) );
  OAI22_X2 U6484 ( .A1(n9447), .A2(n7122), .B1(n12918), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[12]) );
  OAI22_X2 U6485 ( .A1(n9439), .A2(n7147), .B1(n12957), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[5]) );
  OAI22_X2 U6486 ( .A1(n7061), .A2(n7120), .B1(n12933), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[9]) );
  OAI22_X2 U6487 ( .A1(n9338), .A2(n7104), .B1(n9846), .B2(n9391), .ZN(
        pipeline_rs1_data_bypassed[7]) );
  INV_X4 U6488 ( .A(n6636), .ZN(n6637) );
  OAI22_X2 U6489 ( .A1(n9447), .A2(n7145), .B1(n9846), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[7]) );
  INV_X4 U6490 ( .A(n9340), .ZN(imem_haddr[6]) );
  INV_X4 U6491 ( .A(n9344), .ZN(imem_haddr[7]) );
  INV_X4 U6492 ( .A(n9356), .ZN(imem_haddr[11]) );
  INV_X4 U6493 ( .A(n9352), .ZN(imem_haddr[13]) );
  INV_X4 U6494 ( .A(n9350), .ZN(imem_haddr[14]) );
  INV_X4 U6495 ( .A(n9346), .ZN(imem_haddr[16]) );
  INV_X8 U6496 ( .A(n10808), .ZN(imem_haddr[17]) );
  INV_X4 U6497 ( .A(n6956), .ZN(n5963) );
  AOI22_X2 U6498 ( .A1(pipeline_PC_IF_8_), .A2(n9495), .B1(n6737), .B2(
        imem_haddr[8]), .ZN(n6956) );
  INV_X4 U6499 ( .A(n6570), .ZN(n11510) );
  NOR2_X1 U6500 ( .A1(n12501), .A2(n9485), .ZN(n12502) );
  INV_X4 U6501 ( .A(pipeline_rs1_data_bypassed[9]), .ZN(n12501) );
  NOR2_X1 U6502 ( .A1(n12526), .A2(n9486), .ZN(n12527) );
  OAI22_X2 U6503 ( .A1(n718), .A2(n9445), .B1(n12526), .B2(n9785), .ZN(
        pipeline_alu_src_a[3]) );
  AND4_X4 U6504 ( .A1(n7345), .A2(n7346), .A3(n7347), .A4(n7348), .ZN(n7071)
         );
  NOR2_X1 U6505 ( .A1(n12422), .A2(n9484), .ZN(n12423) );
  AOI221_X2 U6506 ( .B1(pipeline_PC_DX[21]), .B2(n9480), .C1(
        pipeline_handler_PC[21]), .C2(n6630), .A(n12455), .ZN(n12456) );
  NAND2_X2 U6507 ( .A1(n6623), .A2(n9486), .ZN(n12554) );
  NOR2_X1 U6508 ( .A1(n12430), .A2(n9484), .ZN(n12431) );
  OAI22_X2 U6509 ( .A1(n719), .A2(n9445), .B1(n12522), .B2(n9785), .ZN(
        pipeline_alu_src_a[4]) );
  AND4_X2 U6510 ( .A1(n7665), .A2(n7666), .A3(n7667), .A4(n7668), .ZN(n7095)
         );
  AOI221_X1 U6511 ( .B1(pipeline_regfile_data[942]), .B2(n6728), .C1(
        pipeline_regfile_data[686]), .C2(n6720), .A(n7669), .ZN(n7668) );
  AND2_X2 U6512 ( .A1(n8379), .A2(n8380), .ZN(n8378) );
  NAND2_X1 U6513 ( .A1(n9489), .A2(pipeline_alu_src_a[9]), .ZN(n11719) );
  NOR2_X1 U6514 ( .A1(pipeline_rs1_data_bypassed[9]), .A2(n9463), .ZN(n10580)
         );
  OAI22_X2 U6515 ( .A1(n10057), .A2(n10242), .B1(n12686), .B2(n10056), .ZN(
        n13159) );
  OAI22_X2 U6516 ( .A1(n9916), .A2(n10056), .B1(n713), .B2(n9915), .ZN(
        pipeline_alu_src_b[10]) );
  AOI221_X1 U6517 ( .B1(pipeline_regfile_data[328]), .B2(n9324), .C1(
        pipeline_regfile_data[264]), .C2(n9327), .A(n8541), .ZN(n8536) );
  AOI221_X1 U6518 ( .B1(pipeline_regfile_data[330]), .B2(n9324), .C1(
        pipeline_regfile_data[266]), .C2(n9327), .A(n8605), .ZN(n8600) );
  INV_X4 U6519 ( .A(pipeline_alu_src_a[5]), .ZN(n6619) );
  INV_X1 U6520 ( .A(n6619), .ZN(n6620) );
  INV_X1 U6521 ( .A(n6619), .ZN(n6621) );
  NAND3_X2 U6522 ( .A1(pipeline_regfile_N17), .A2(pipeline_regfile_N19), .A3(
        n6628), .ZN(n8232) );
  AND2_X1 U6523 ( .A1(pipeline_regfile_N17), .A2(pipeline_regfile_N18), .ZN(
        n7175) );
  INV_X8 U6524 ( .A(n9362), .ZN(imem_haddr[19]) );
  INV_X8 U6525 ( .A(n9366), .ZN(imem_haddr[22]) );
  INV_X8 U6526 ( .A(n9374), .ZN(imem_haddr[18]) );
  INV_X8 U6527 ( .A(n9376), .ZN(imem_haddr[21]) );
  INV_X8 U6528 ( .A(n9368), .ZN(imem_haddr[20]) );
  NAND2_X1 U6529 ( .A1(pipeline_regfile_N18), .A2(n6745), .ZN(n12825) );
  NOR3_X1 U6530 ( .A1(pipeline_ctrl_N81), .A2(pipeline_regfile_N18), .A3(
        pipeline_ctrl_N82), .ZN(n9621) );
  NAND2_X1 U6531 ( .A1(n9790), .A2(pipeline_regfile_N18), .ZN(n9715) );
  AND2_X4 U6532 ( .A1(pipeline_regfile_N18), .A2(n702), .ZN(n7174) );
  INV_X4 U6533 ( .A(n9398), .ZN(n9399) );
  AOI22_X2 U6534 ( .A1(n6927), .A2(n9458), .B1(pipeline_alu_src_b[4]), .B2(
        n9452), .ZN(n9388) );
  AOI221_X2 U6535 ( .B1(pipeline_regfile_data[955]), .B2(n6728), .C1(
        pipeline_regfile_data[699]), .C2(n6720), .A(n8083), .ZN(n8082) );
  NAND2_X2 U6536 ( .A1(n7170), .A2(pipeline_regfile_N14), .ZN(n9294) );
  INV_X1 U6537 ( .A(n9481), .ZN(n6622) );
  INV_X2 U6538 ( .A(n6556), .ZN(n12299) );
  AND4_X2 U6539 ( .A1(n7473), .A2(n7474), .A3(n7475), .A4(n7476), .ZN(n7139)
         );
  AOI221_X2 U6540 ( .B1(pipeline_regfile_data[355]), .B2(n8249), .C1(
        pipeline_regfile_data[291]), .C2(n8253), .A(n7322), .ZN(n7321) );
  AND4_X2 U6541 ( .A1(n8079), .A2(n8080), .A3(n8081), .A4(n8082), .ZN(n7125)
         );
  INV_X2 U6542 ( .A(n6622), .ZN(n6623) );
  AND2_X2 U6543 ( .A1(n8315), .A2(n8316), .ZN(n8314) );
  INV_X4 U6544 ( .A(pipeline_alu_src_a[22]), .ZN(n6624) );
  INV_X1 U6545 ( .A(n6624), .ZN(n6625) );
  INV_X1 U6546 ( .A(n6624), .ZN(n6626) );
  AND4_X2 U6547 ( .A1(n7281), .A2(n7282), .A3(n7283), .A4(n7284), .ZN(n7096)
         );
  OAI22_X2 U6548 ( .A1(n9859), .A2(n10056), .B1(n9632), .B2(n9915), .ZN(
        pipeline_alu_src_b[9]) );
  INV_X2 U6549 ( .A(n13159), .ZN(n12566) );
  INV_X2 U6550 ( .A(n700), .ZN(n6627) );
  INV_X4 U6551 ( .A(n6627), .ZN(n6628) );
  AOI221_X1 U6552 ( .B1(pipeline_md_N38), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[9]), .A(n10556), .ZN(n10557) );
  AOI221_X2 U6553 ( .B1(n9483), .B2(n6637), .C1(pipeline_PC_DX[1]), .C2(n9480), 
        .A(n12536), .ZN(n12537) );
  NAND2_X1 U6554 ( .A1(n9483), .A2(pipeline_imm_31_), .ZN(n12553) );
  NAND2_X1 U6555 ( .A1(n12588), .A2(n13159), .ZN(n12589) );
  OAI22_X2 U6556 ( .A1(n9439), .A2(n7091), .B1(n9825), .B2(n9392), .ZN(
        pipeline_rs1_data_bypassed[16]) );
  NOR2_X1 U6557 ( .A1(pipeline_rs1_data_bypassed[15]), .A2(n9463), .ZN(n11122)
         );
  AOI221_X1 U6558 ( .B1(pipeline_md_N44), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[15]), .A(n11096), .ZN(n11097) );
  OAI22_X1 U6559 ( .A1(n9338), .A2(n7097), .B1(n12977), .B2(n9391), .ZN(
        pipeline_rs1_data_bypassed[1]) );
  OAI22_X1 U6560 ( .A1(n9338), .A2(n7106), .B1(n9954), .B2(n9392), .ZN(
        pipeline_rs1_data_bypassed[18]) );
  OAI22_X1 U6561 ( .A1(n9338), .A2(n7112), .B1(n9985), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[22]) );
  NAND3_X1 U6562 ( .A1(n637), .A2(n636), .A3(n9614), .ZN(n10258) );
  NOR2_X2 U6563 ( .A1(n12485), .A2(n9485), .ZN(n12486) );
  NOR2_X1 U6564 ( .A1(n700), .A2(n702), .ZN(n6940) );
  AND3_X1 U6565 ( .A1(n6628), .A2(n10336), .A3(n6796), .ZN(n7193) );
  OAI22_X1 U6566 ( .A1(n6628), .A2(n12562), .B1(n595), .B2(n12561), .ZN(
        pipeline_PCmux_offset[1]) );
  INV_X8 U6567 ( .A(n12532), .ZN(n6629) );
  INV_X16 U6568 ( .A(n6629), .ZN(n6630) );
  INV_X2 U6569 ( .A(n12410), .ZN(n12532) );
  OAI221_X2 U6570 ( .B1(n9487), .B2(n12488), .C1(n1496), .C2(n6661), .A(n12487), .ZN(pipeline_PCmux_base[13]) );
  AOI221_X1 U6571 ( .B1(pipeline_md_N36), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[7]), .A(n10665), .ZN(n10666) );
  NOR2_X1 U6572 ( .A1(pipeline_rs1_data_bypassed[7]), .A2(n9463), .ZN(n10688)
         );
  INV_X1 U6573 ( .A(n6631), .ZN(n6632) );
  NOR2_X1 U6574 ( .A1(pipeline_alu_src_b[22]), .A2(n12357), .ZN(n11762) );
  NAND3_X2 U6575 ( .A1(n9885), .A2(n9886), .A3(n9884), .ZN(n9898) );
  AOI221_X1 U6576 ( .B1(pipeline_regfile_data[113]), .B2(n8247), .C1(
        pipeline_regfile_data[49]), .C2(n8253), .A(n7777), .ZN(n7776) );
  AOI221_X1 U6577 ( .B1(pipeline_regfile_data[369]), .B2(n8247), .C1(
        pipeline_regfile_data[305]), .C2(n8253), .A(n7769), .ZN(n7768) );
  AOI221_X1 U6578 ( .B1(pipeline_regfile_data[111]), .B2(n8247), .C1(
        pipeline_regfile_data[47]), .C2(n8253), .A(n7714), .ZN(n7713) );
  AOI221_X1 U6579 ( .B1(pipeline_regfile_data[106]), .B2(n8248), .C1(
        pipeline_regfile_data[42]), .C2(n8253), .A(n7554), .ZN(n7553) );
  AOI221_X1 U6580 ( .B1(pipeline_regfile_data[361]), .B2(n8248), .C1(
        pipeline_regfile_data[297]), .C2(n8253), .A(n7514), .ZN(n7513) );
  AOI221_X1 U6581 ( .B1(pipeline_regfile_data[103]), .B2(n8248), .C1(
        pipeline_regfile_data[39]), .C2(n8253), .A(n7458), .ZN(n7457) );
  AOI221_X1 U6582 ( .B1(pipeline_regfile_data[101]), .B2(n8249), .C1(
        pipeline_regfile_data[37]), .C2(n8253), .A(n7394), .ZN(n7393) );
  AOI221_X1 U6583 ( .B1(pipeline_regfile_data[104]), .B2(n8248), .C1(
        pipeline_regfile_data[40]), .C2(n8253), .A(n7490), .ZN(n7489) );
  AOI221_X1 U6584 ( .B1(pipeline_regfile_data[366]), .B2(n8247), .C1(
        pipeline_regfile_data[302]), .C2(n8253), .A(n7674), .ZN(n7673) );
  AOI221_X1 U6585 ( .B1(pipeline_regfile_data[357]), .B2(n8249), .C1(
        pipeline_regfile_data[293]), .C2(n8253), .A(n7386), .ZN(n7385) );
  AOI221_X1 U6586 ( .B1(pipeline_regfile_data[360]), .B2(n8248), .C1(
        pipeline_regfile_data[296]), .C2(n8253), .A(n7482), .ZN(n7481) );
  AND4_X2 U6587 ( .A1(n8401), .A2(n8402), .A3(n8403), .A4(n8404), .ZN(n7070)
         );
  INV_X4 U6588 ( .A(pipeline_alu_src_a[3]), .ZN(n6633) );
  INV_X1 U6589 ( .A(n6633), .ZN(n6634) );
  INV_X1 U6590 ( .A(n6633), .ZN(n6635) );
  INV_X4 U6591 ( .A(pipeline_rs1_data_bypassed[1]), .ZN(n6636) );
  AOI221_X1 U6592 ( .B1(pipeline_regfile_data[87]), .B2(n9323), .C1(
        pipeline_regfile_data[23]), .C2(n9326), .A(n9027), .ZN(n9022) );
  AOI221_X1 U6593 ( .B1(pipeline_regfile_data[90]), .B2(n9324), .C1(
        pipeline_regfile_data[26]), .C2(n9327), .A(n9123), .ZN(n9118) );
  AOI221_X1 U6594 ( .B1(pipeline_regfile_data[86]), .B2(n9323), .C1(
        pipeline_regfile_data[22]), .C2(n9327), .A(n8995), .ZN(n8990) );
  AOI221_X1 U6595 ( .B1(pipeline_regfile_data[119]), .B2(n9308), .C1(
        pipeline_regfile_data[55]), .C2(n9314), .A(n9024), .ZN(n9023) );
  AOI221_X1 U6596 ( .B1(pipeline_regfile_data[375]), .B2(n9308), .C1(
        pipeline_regfile_data[311]), .C2(n9314), .A(n9016), .ZN(n9015) );
  AOI221_X1 U6597 ( .B1(pipeline_regfile_data[118]), .B2(n9308), .C1(
        pipeline_regfile_data[54]), .C2(n9314), .A(n8992), .ZN(n8991) );
  AOI221_X1 U6598 ( .B1(pipeline_regfile_data[374]), .B2(n9308), .C1(
        pipeline_regfile_data[310]), .C2(n9314), .A(n8984), .ZN(n8983) );
  AOI221_X1 U6599 ( .B1(pipeline_regfile_data[121]), .B2(n9308), .C1(
        pipeline_regfile_data[57]), .C2(n9314), .A(n9088), .ZN(n9087) );
  AOI221_X1 U6600 ( .B1(pipeline_regfile_data[120]), .B2(n9308), .C1(
        pipeline_regfile_data[56]), .C2(n9314), .A(n9056), .ZN(n9055) );
  AOI221_X1 U6601 ( .B1(pipeline_regfile_data[377]), .B2(n9308), .C1(
        pipeline_regfile_data[313]), .C2(n9314), .A(n9080), .ZN(n9079) );
  AOI221_X1 U6602 ( .B1(pipeline_regfile_data[116]), .B2(n9308), .C1(
        pipeline_regfile_data[52]), .C2(n9314), .A(n8930), .ZN(n8929) );
  AOI221_X1 U6603 ( .B1(pipeline_regfile_data[117]), .B2(n9308), .C1(
        pipeline_regfile_data[53]), .C2(n9314), .A(n8962), .ZN(n8961) );
  AOI221_X1 U6604 ( .B1(pipeline_regfile_data[373]), .B2(n9308), .C1(
        pipeline_regfile_data[309]), .C2(n9314), .A(n8954), .ZN(n8953) );
  AOI221_X1 U6605 ( .B1(pipeline_regfile_data[115]), .B2(n9308), .C1(
        pipeline_regfile_data[51]), .C2(n9314), .A(n8898), .ZN(n8897) );
  AOI221_X1 U6606 ( .B1(pipeline_regfile_data[376]), .B2(n9308), .C1(
        pipeline_regfile_data[312]), .C2(n9314), .A(n9048), .ZN(n9047) );
  AOI221_X1 U6607 ( .B1(pipeline_regfile_data[367]), .B2(n9309), .C1(
        pipeline_regfile_data[303]), .C2(n9314), .A(n8762), .ZN(n8761) );
  NAND2_X2 U6608 ( .A1(n6575), .A2(n9723), .ZN(n6638) );
  NAND2_X4 U6609 ( .A1(n6575), .A2(n9723), .ZN(n10055) );
  NAND2_X2 U6610 ( .A1(n10098), .A2(n12832), .ZN(n6639) );
  INV_X4 U6611 ( .A(n9294), .ZN(n9318) );
  AND3_X4 U6612 ( .A1(n7051), .A2(n10251), .A3(n9402), .ZN(n6640) );
  AND3_X4 U6613 ( .A1(n713), .A2(n10242), .A3(n7055), .ZN(n6641) );
  NAND3_X1 U6614 ( .A1(pipeline_regfile_N18), .A2(n702), .A3(n693), .ZN(n6642)
         );
  AND2_X4 U6615 ( .A1(n9518), .A2(n12828), .ZN(n6643) );
  AND2_X4 U6616 ( .A1(n6716), .A2(n6852), .ZN(n6644) );
  AND2_X4 U6617 ( .A1(n6716), .A2(n6853), .ZN(n6645) );
  AND2_X4 U6618 ( .A1(n6716), .A2(n6856), .ZN(n6646) );
  AND2_X4 U6619 ( .A1(n6716), .A2(n6859), .ZN(n6647) );
  AND2_X4 U6620 ( .A1(n6716), .A2(n6855), .ZN(n6648) );
  AND2_X4 U6621 ( .A1(n6852), .A2(n6717), .ZN(n6649) );
  AND2_X4 U6622 ( .A1(n6853), .A2(n6717), .ZN(n6650) );
  AND2_X4 U6623 ( .A1(n6856), .A2(n6717), .ZN(n6651) );
  AND2_X4 U6624 ( .A1(n6859), .A2(n6717), .ZN(n6652) );
  AND2_X4 U6625 ( .A1(n6716), .A2(n6854), .ZN(n6653) );
  AND2_X4 U6626 ( .A1(n6855), .A2(n6717), .ZN(n6654) );
  AND2_X4 U6627 ( .A1(n6854), .A2(n6717), .ZN(n6655) );
  AND2_X4 U6628 ( .A1(n6716), .A2(n6756), .ZN(n6656) );
  AND2_X4 U6629 ( .A1(n6716), .A2(n6757), .ZN(n6657) );
  AND2_X4 U6630 ( .A1(n6756), .A2(n6717), .ZN(n6658) );
  NAND2_X4 U6631 ( .A1(n6753), .A2(n6689), .ZN(n6659) );
  NAND2_X4 U6632 ( .A1(n9516), .A2(n13130), .ZN(n6660) );
  NAND2_X4 U6633 ( .A1(n12412), .A2(n12560), .ZN(n6661) );
  NAND2_X4 U6634 ( .A1(n10388), .A2(n13130), .ZN(n6662) );
  NAND2_X4 U6635 ( .A1(pipeline_regfile_N20), .A2(n8214), .ZN(n6663) );
  INV_X4 U6636 ( .A(n9317), .ZN(n9320) );
  AND2_X4 U6637 ( .A1(pipeline_inst_DX[25]), .A2(n6711), .ZN(n6664) );
  AND2_X4 U6638 ( .A1(n7168), .A2(n3704), .ZN(n6665) );
  AND2_X4 U6639 ( .A1(n6698), .A2(n603), .ZN(n6666) );
  NAND2_X4 U6640 ( .A1(n10271), .A2(n10277), .ZN(n6667) );
  NOR2_X4 U6641 ( .A1(n11285), .A2(n11199), .ZN(n6668) );
  NOR2_X4 U6642 ( .A1(n11200), .A2(n11199), .ZN(n6669) );
  AND3_X4 U6643 ( .A1(n11193), .A2(n12806), .A3(n9515), .ZN(n6670) );
  AND2_X4 U6644 ( .A1(n7088), .A2(n6855), .ZN(n6671) );
  AND2_X4 U6645 ( .A1(n7088), .A2(n6756), .ZN(n6672) );
  AND2_X4 U6646 ( .A1(n7087), .A2(n6852), .ZN(n6673) );
  AND2_X4 U6647 ( .A1(n7087), .A2(n6853), .ZN(n6674) );
  AND2_X4 U6648 ( .A1(n7087), .A2(n6856), .ZN(n6675) );
  AND2_X4 U6649 ( .A1(n7087), .A2(n6859), .ZN(n6676) );
  AND2_X4 U6650 ( .A1(n7087), .A2(n6855), .ZN(n6677) );
  AND2_X4 U6651 ( .A1(n7087), .A2(n6854), .ZN(n6678) );
  AND2_X4 U6652 ( .A1(n7087), .A2(n6756), .ZN(n6679) );
  AND2_X4 U6653 ( .A1(n7087), .A2(n6757), .ZN(n6680) );
  AND2_X4 U6654 ( .A1(n7088), .A2(n6852), .ZN(n6681) );
  AND2_X4 U6655 ( .A1(n7088), .A2(n6853), .ZN(n6682) );
  AND2_X4 U6656 ( .A1(n7088), .A2(n6856), .ZN(n6683) );
  AND2_X4 U6657 ( .A1(n7088), .A2(n6859), .ZN(n6684) );
  AND2_X4 U6658 ( .A1(n7088), .A2(n6854), .ZN(n6685) );
  AND2_X4 U6659 ( .A1(n7088), .A2(n6757), .ZN(n6686) );
  NAND2_X4 U6660 ( .A1(n6799), .A2(n6705), .ZN(n6687) );
  NAND2_X4 U6661 ( .A1(n9530), .A2(n13130), .ZN(n6688) );
  NAND2_X4 U6662 ( .A1(n6753), .A2(n10825), .ZN(n6689) );
  NAND2_X4 U6663 ( .A1(n6708), .A2(n13130), .ZN(n6690) );
  NAND2_X4 U6664 ( .A1(n9523), .A2(n8223), .ZN(n6691) );
  NAND2_X4 U6665 ( .A1(n6914), .A2(n10270), .ZN(n6692) );
  NAND2_X4 U6666 ( .A1(n9500), .A2(n6917), .ZN(n6693) );
  NAND2_X4 U6667 ( .A1(n784), .A2(n9534), .ZN(n6694) );
  NAND2_X4 U6668 ( .A1(n8223), .A2(n8214), .ZN(n6695) );
  INV_X4 U6669 ( .A(n9307), .ZN(n9308) );
  INV_X4 U6670 ( .A(n12556), .ZN(n9483) );
  NAND2_X2 U6671 ( .A1(pipeline_regfile_N17), .A2(n6940), .ZN(n6696) );
  AND2_X4 U6672 ( .A1(n7081), .A2(n7169), .ZN(n6697) );
  AND2_X4 U6673 ( .A1(n10260), .A2(n3704), .ZN(n6698) );
  NAND2_X4 U6674 ( .A1(n10278), .A2(n10277), .ZN(n6699) );
  AND2_X4 U6675 ( .A1(n6820), .A2(n6749), .ZN(n6700) );
  AND4_X4 U6676 ( .A1(n10501), .A2(n10500), .A3(n10499), .A4(n10498), .ZN(
        n6701) );
  NAND2_X4 U6677 ( .A1(n9529), .A2(n13130), .ZN(n6702) );
  NAND2_X4 U6678 ( .A1(n3683), .A2(n13130), .ZN(n6703) );
  NAND2_X4 U6679 ( .A1(n10352), .A2(n10522), .ZN(n6704) );
  NAND2_X4 U6680 ( .A1(n6748), .A2(n7165), .ZN(n6705) );
  AND2_X4 U6681 ( .A1(n10777), .A2(n13130), .ZN(n6706) );
  NAND3_X4 U6682 ( .A1(n13139), .A2(n9533), .A3(htif_pcr_req_addr[0]), .ZN(
        n6707) );
  NAND2_X4 U6683 ( .A1(n10263), .A2(n13130), .ZN(n6708) );
  NAND3_X1 U6684 ( .A1(n7193), .A2(n693), .A3(n9402), .ZN(n12258) );
  AND2_X4 U6685 ( .A1(n9326), .A2(n6736), .ZN(n6709) );
  INV_X4 U6686 ( .A(n6779), .ZN(n9447) );
  INV_X4 U6687 ( .A(n6779), .ZN(n7061) );
  NAND2_X1 U6688 ( .A1(n7175), .A2(n702), .ZN(n8240) );
  INV_X4 U6689 ( .A(n7015), .ZN(n8262) );
  AND2_X4 U6690 ( .A1(n10236), .A2(n10338), .ZN(n6711) );
  INV_X4 U6691 ( .A(n6642), .ZN(n8261) );
  INV_X4 U6692 ( .A(n9481), .ZN(n9480) );
  AND2_X4 U6693 ( .A1(n6739), .A2(n7177), .ZN(n6712) );
  AND4_X4 U6694 ( .A1(n11244), .A2(n11243), .A3(n11242), .A4(n11241), .ZN(
        n6713) );
  AND3_X4 U6695 ( .A1(n9469), .A2(n12255), .A3(n6819), .ZN(n6714) );
  OR2_X4 U6696 ( .A1(n6747), .A2(pipeline_md_N21), .ZN(n6715) );
  AND2_X4 U6697 ( .A1(n7191), .A2(n12995), .ZN(n6716) );
  AND2_X4 U6698 ( .A1(n7191), .A2(n12996), .ZN(n6717) );
  AND2_X4 U6699 ( .A1(n8264), .A2(n6774), .ZN(n6719) );
  AND2_X4 U6700 ( .A1(n8257), .A2(n6774), .ZN(n6720) );
  AND2_X4 U6701 ( .A1(n8255), .A2(n6774), .ZN(n6721) );
  AND2_X4 U6702 ( .A1(n8251), .A2(n6775), .ZN(n6722) );
  AND2_X4 U6703 ( .A1(n6599), .A2(n6775), .ZN(n6723) );
  AND2_X4 U6704 ( .A1(n6774), .A2(n8261), .ZN(n6724) );
  AND2_X4 U6705 ( .A1(n8255), .A2(n6775), .ZN(n6725) );
  AND2_X4 U6706 ( .A1(n8253), .A2(n6774), .ZN(n6726) );
  AND2_X4 U6707 ( .A1(n8262), .A2(n6775), .ZN(n6727) );
  AND2_X4 U6708 ( .A1(n8257), .A2(n6775), .ZN(n6728) );
  AND2_X4 U6709 ( .A1(n8261), .A2(n6775), .ZN(n6729) );
  AND2_X4 U6710 ( .A1(n8245), .A2(n6774), .ZN(n6730) );
  AND2_X4 U6711 ( .A1(n8269), .A2(n6774), .ZN(n6731) );
  AND2_X4 U6712 ( .A1(n8245), .A2(n6775), .ZN(n6732) );
  AND2_X4 U6713 ( .A1(n8271), .A2(n6775), .ZN(n6733) );
  AND2_X4 U6714 ( .A1(n6599), .A2(n6774), .ZN(n6734) );
  AND2_X4 U6715 ( .A1(n7077), .A2(n9402), .ZN(n6735) );
  AND2_X4 U6716 ( .A1(pipeline_regfile_N16), .A2(n9279), .ZN(n6736) );
  AND2_X4 U6717 ( .A1(n10386), .A2(n13130), .ZN(n6737) );
  INV_X4 U6718 ( .A(n6776), .ZN(n9306) );
  INV_X4 U6719 ( .A(n8240), .ZN(n8245) );
  AND2_X4 U6720 ( .A1(pipeline_dmem_type_2_), .A2(dmem_hsize[1]), .ZN(n6738)
         );
  AND2_X4 U6721 ( .A1(n9628), .A2(n12834), .ZN(n6739) );
  INV_X4 U6722 ( .A(n9313), .ZN(n9312) );
  AND4_X4 U6723 ( .A1(n9652), .A2(n9670), .A3(n10131), .A4(n6739), .ZN(n6740)
         );
  NAND2_X1 U6724 ( .A1(n7170), .A2(n638), .ZN(n9298) );
  AND2_X4 U6725 ( .A1(n6784), .A2(pipeline_inst_DX[30]), .ZN(n6741) );
  INV_X4 U6726 ( .A(n13182), .ZN(n9360) );
  AND2_X4 U6727 ( .A1(n6799), .A2(n12404), .ZN(n6742) );
  AND2_X4 U6728 ( .A1(n10127), .A2(n6799), .ZN(n6743) );
  NAND3_X2 U6729 ( .A1(n9801), .A2(n6578), .A3(n9800), .ZN(n6744) );
  AND4_X4 U6730 ( .A1(n6794), .A2(n13096), .A3(n9618), .A4(n10132), .ZN(n6745)
         );
  AND2_X4 U6731 ( .A1(n11578), .A2(n11641), .ZN(n6746) );
  AND3_X4 U6732 ( .A1(n3785), .A2(n8223), .A3(n7166), .ZN(n6748) );
  AND2_X4 U6733 ( .A1(n10350), .A2(n10353), .ZN(n6749) );
  AND2_X4 U6734 ( .A1(n6687), .A2(n6705), .ZN(n6750) );
  AND2_X4 U6735 ( .A1(n4184), .A2(n13130), .ZN(n6753) );
  AND2_X4 U6736 ( .A1(n6916), .A2(n10275), .ZN(n6754) );
  AND2_X4 U6737 ( .A1(n6916), .A2(n10270), .ZN(n6755) );
  AND2_X4 U6738 ( .A1(n6912), .A2(n12990), .ZN(n6756) );
  AND2_X4 U6739 ( .A1(n6912), .A2(n12991), .ZN(n6757) );
  AND2_X4 U6740 ( .A1(n9320), .A2(n6736), .ZN(n6761) );
  AND2_X4 U6741 ( .A1(n6736), .A2(n9325), .ZN(n6762) );
  AND2_X4 U6742 ( .A1(n9328), .A2(n7164), .ZN(n6763) );
  AND2_X4 U6743 ( .A1(n9321), .A2(n6736), .ZN(n6764) );
  AND2_X4 U6744 ( .A1(n9319), .A2(n7164), .ZN(n6765) );
  AND2_X4 U6745 ( .A1(n9327), .A2(n7164), .ZN(n6766) );
  AND2_X4 U6746 ( .A1(n9321), .A2(n7164), .ZN(n6767) );
  OAI22_X2 U6747 ( .A1(n724), .A2(n9445), .B1(n12501), .B2(n9443), .ZN(
        pipeline_alu_src_a[9]) );
  AND2_X4 U6748 ( .A1(n9324), .A2(n7164), .ZN(n6768) );
  AND2_X4 U6749 ( .A1(n9331), .A2(n6736), .ZN(n6769) );
  AND2_X4 U6750 ( .A1(n9309), .A2(n7164), .ZN(n6770) );
  OAI22_X2 U6751 ( .A1(n9855), .A2(n9448), .B1(n9634), .B2(n9915), .ZN(
        pipeline_alu_src_b[8]) );
  AND2_X4 U6752 ( .A1(n9330), .A2(n7164), .ZN(n6772) );
  AND2_X4 U6753 ( .A1(n9328), .A2(n6736), .ZN(n6773) );
  INV_X4 U6754 ( .A(n13160), .ZN(n12563) );
  AND2_X4 U6755 ( .A1(pipeline_regfile_N21), .A2(n8223), .ZN(n6774) );
  AND2_X4 U6756 ( .A1(pipeline_regfile_N21), .A2(pipeline_regfile_N20), .ZN(
        n6775) );
  AND2_X4 U6757 ( .A1(pipeline_regfile_N15), .A2(n9270), .ZN(n6776) );
  AND2_X4 U6758 ( .A1(n12832), .A2(n6662), .ZN(n6777) );
  NAND2_X2 U6759 ( .A1(n9459), .A2(pipeline_alu_src_a[0]), .ZN(n6778) );
  AND2_X4 U6760 ( .A1(n6638), .A2(n9703), .ZN(n6779) );
  AND2_X4 U6761 ( .A1(n12408), .A2(n12407), .ZN(n6780) );
  OAI22_X2 U6762 ( .A1(n11809), .A2(n9455), .B1(n6604), .B2(n9451), .ZN(n9899)
         );
  AND2_X4 U6763 ( .A1(n12554), .A2(pipeline_imm_31_), .ZN(n6781) );
  OR3_X2 U6764 ( .A1(n6993), .A2(n6994), .A3(n8312), .ZN(n6782) );
  OR3_X4 U6765 ( .A1(n7010), .A2(n7011), .A3(n8051), .ZN(n6783) );
  AND3_X4 U6766 ( .A1(pipeline_dmem_type_2_), .A2(n602), .A3(dmem_hsize[0]), 
        .ZN(n6784) );
  NAND3_X2 U6767 ( .A1(n6999), .A2(n7000), .A3(n7001), .ZN(n6785) );
  OR2_X4 U6768 ( .A1(n9582), .A2(n9583), .ZN(n6786) );
  INV_X4 U6769 ( .A(n9887), .ZN(n9885) );
  AND4_X4 U6770 ( .A1(n8561), .A2(n8562), .A3(n8563), .A4(n8564), .ZN(n6787)
         );
  AND4_X4 U6771 ( .A1(n9135), .A2(n9136), .A3(n9137), .A4(n9138), .ZN(n6788)
         );
  AND4_X4 U6772 ( .A1(n7217), .A2(n7218), .A3(n7219), .A4(n7220), .ZN(n6789)
         );
  AND4_X4 U6773 ( .A1(n8372), .A2(n8373), .A3(n8374), .A4(n8375), .ZN(n6790)
         );
  INV_X4 U6774 ( .A(n7053), .ZN(n9313) );
  AND2_X4 U6775 ( .A1(n9895), .A2(n9896), .ZN(n6791) );
  NAND2_X2 U6776 ( .A1(n7052), .A2(n9722), .ZN(n6792) );
  INV_X4 U6777 ( .A(n6696), .ZN(n8254) );
  AND2_X4 U6778 ( .A1(n6665), .A2(pipeline_dmem_type_2_), .ZN(n6793) );
  OAI22_X2 U6779 ( .A1(n7061), .A2(n7130), .B1(n9819), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[17]) );
  AND4_X4 U6780 ( .A1(n595), .A2(n594), .A3(n596), .A4(n9615), .ZN(n6794) );
  AND2_X4 U6781 ( .A1(dmem_hsize[1]), .A2(n603), .ZN(n6795) );
  AND2_X4 U6782 ( .A1(n10337), .A2(n10338), .ZN(n6796) );
  AND2_X4 U6783 ( .A1(n12684), .A2(n13034), .ZN(n6797) );
  AND3_X4 U6784 ( .A1(n10264), .A2(n7183), .A3(n9504), .ZN(n6798) );
  AND2_X4 U6785 ( .A1(n12149), .A2(n6369), .ZN(n6799) );
  AND4_X4 U6786 ( .A1(n11777), .A2(n11776), .A3(n11775), .A4(n11774), .ZN(
        n6800) );
  AND4_X4 U6787 ( .A1(n11718), .A2(n11717), .A3(n11716), .A4(n11715), .ZN(
        n6801) );
  AND2_X4 U6788 ( .A1(n12020), .A2(n12026), .ZN(n6802) );
  AND2_X4 U6789 ( .A1(n12795), .A2(n11772), .ZN(n6803) );
  AND4_X4 U6790 ( .A1(n11961), .A2(n11960), .A3(n11959), .A4(n11958), .ZN(
        n6804) );
  AND4_X4 U6791 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n6805) );
  AND2_X4 U6792 ( .A1(n11503), .A2(n11502), .ZN(n6806) );
  AND2_X4 U6793 ( .A1(n10184), .A2(n9620), .ZN(n6807) );
  AND3_X4 U6794 ( .A1(n7183), .A2(n10265), .A3(n9504), .ZN(n6808) );
  AND2_X4 U6795 ( .A1(n10277), .A2(n10201), .ZN(n6809) );
  AND4_X4 U6796 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(
        n6811) );
  AND2_X4 U6797 ( .A1(n7069), .A2(n10083), .ZN(n6812) );
  AND2_X4 U6798 ( .A1(n7069), .A2(n10085), .ZN(n6813) );
  OR2_X4 U6799 ( .A1(n6747), .A2(n13128), .ZN(n6814) );
  AND4_X4 U6800 ( .A1(n10790), .A2(n10789), .A3(n10788), .A4(n10787), .ZN(
        n6816) );
  AND2_X4 U6801 ( .A1(n7063), .A2(n11111), .ZN(n6818) );
  AND2_X4 U6802 ( .A1(n10419), .A2(n12612), .ZN(n6819) );
  AND2_X4 U6803 ( .A1(n10335), .A2(n9492), .ZN(n6820) );
  AND2_X4 U6804 ( .A1(n11321), .A2(n11320), .ZN(n6821) );
  AND2_X4 U6805 ( .A1(n6748), .A2(n7169), .ZN(n6826) );
  AND2_X4 U6806 ( .A1(n10824), .A2(n6641), .ZN(n6843) );
  AND3_X4 U6807 ( .A1(n799), .A2(n7083), .A3(n9525), .ZN(n6844) );
  AND2_X4 U6808 ( .A1(n10824), .A2(n7193), .ZN(n6847) );
  AND2_X4 U6809 ( .A1(n12905), .A2(n12981), .ZN(n6848) );
  AND4_X4 U6810 ( .A1(n3785), .A2(n13130), .A3(n6697), .A4(n8223), .ZN(n6849)
         );
  AND3_X4 U6811 ( .A1(pipeline_reg_to_wr_WB[1]), .A2(n12990), .A3(
        pipeline_reg_to_wr_WB[2]), .ZN(n6852) );
  AND3_X4 U6812 ( .A1(pipeline_reg_to_wr_WB[1]), .A2(n12991), .A3(
        pipeline_reg_to_wr_WB[2]), .ZN(n6853) );
  AND3_X4 U6813 ( .A1(pipeline_reg_to_wr_WB[1]), .A2(n12988), .A3(n12991), 
        .ZN(n6854) );
  AND3_X4 U6814 ( .A1(n12988), .A2(n12990), .A3(pipeline_reg_to_wr_WB[1]), 
        .ZN(n6855) );
  AND3_X4 U6815 ( .A1(n12989), .A2(n12990), .A3(pipeline_reg_to_wr_WB[2]), 
        .ZN(n6856) );
  AND3_X4 U6816 ( .A1(n12989), .A2(n12991), .A3(pipeline_reg_to_wr_WB[2]), 
        .ZN(n6859) );
  AND2_X4 U6817 ( .A1(n12989), .A2(n12988), .ZN(n6912) );
  AND2_X4 U6818 ( .A1(n962), .A2(n10269), .ZN(n6914) );
  AND2_X4 U6819 ( .A1(n10192), .A2(n10269), .ZN(n6916) );
  AND2_X4 U6820 ( .A1(n6914), .A2(n10275), .ZN(n6917) );
  AND2_X4 U6821 ( .A1(n10198), .A2(n9519), .ZN(n6918) );
  OAI22_X2 U6822 ( .A1(n12530), .A2(n9785), .B1(n9786), .B2(n717), .ZN(
        pipeline_alu_src_a[2]) );
  AOI22_X2 U6823 ( .A1(pipeline_rs1_data_bypassed[12]), .A2(n9444), .B1(n9446), 
        .B2(pipeline_PC_DX[12]), .ZN(n6924) );
  INV_X4 U6824 ( .A(n6924), .ZN(pipeline_alu_src_a[12]) );
  INV_X4 U6825 ( .A(n9786), .ZN(n9446) );
  INV_X4 U6826 ( .A(pipeline_alu_src_a[20]), .ZN(n6925) );
  AOI22_X2 U6827 ( .A1(pipeline_alu_src_a[12]), .A2(n9457), .B1(
        pipeline_alu_src_b[12]), .B2(n9452), .ZN(n6926) );
  INV_X4 U6828 ( .A(n6926), .ZN(n9934) );
  INV_X4 U6829 ( .A(pipeline_alu_src_b[12]), .ZN(n11656) );
  OAI221_X2 U6830 ( .B1(n9912), .B2(n10056), .C1(n601), .C2(n9396), .A(n9967), 
        .ZN(pipeline_alu_src_b[12]) );
  NAND2_X2 U6831 ( .A1(n9930), .A2(n9929), .ZN(n9938) );
  NAND3_X2 U6832 ( .A1(n7007), .A2(n7008), .A3(n9706), .ZN(n6929) );
  INV_X4 U6833 ( .A(n6929), .ZN(n7009) );
  INV_X4 U6834 ( .A(n6930), .ZN(n8981) );
  NAND2_X2 U6835 ( .A1(n8990), .A2(n8991), .ZN(n6931) );
  NAND2_X2 U6836 ( .A1(n8982), .A2(n8983), .ZN(n6932) );
  INV_X4 U6837 ( .A(n7015), .ZN(n8263) );
  INV_X4 U6838 ( .A(n7015), .ZN(n8265) );
  NAND3_X1 U6839 ( .A1(n702), .A2(n693), .A3(n9658), .ZN(n7015) );
  OAI221_X2 U6840 ( .B1(n6934), .B2(n9293), .C1(n6935), .C2(n9292), .A(n6936), 
        .ZN(n6933) );
  NAND2_X2 U6841 ( .A1(pipeline_regfile_data[611]), .A2(n8302), .ZN(n6936) );
  INV_X4 U6842 ( .A(n9293), .ZN(n8299) );
  NAND2_X2 U6843 ( .A1(n9313), .A2(n6736), .ZN(n9293) );
  INV_X4 U6844 ( .A(n9292), .ZN(n8300) );
  INV_X4 U6845 ( .A(n9333), .ZN(n9330) );
  INV_X4 U6846 ( .A(n7171), .ZN(n9333) );
  INV_X4 U6847 ( .A(n12265), .ZN(n9398) );
  AND2_X2 U6848 ( .A1(n7672), .A2(n7673), .ZN(n7671) );
  INV_X2 U6849 ( .A(n12554), .ZN(n12555) );
  NOR2_X2 U6850 ( .A1(n9875), .A2(n9874), .ZN(n9876) );
  NOR2_X1 U6851 ( .A1(n6937), .A2(n9291), .ZN(n8426) );
  NAND3_X2 U6852 ( .A1(n9885), .A2(n9890), .A3(n9889), .ZN(n9897) );
  NAND2_X2 U6853 ( .A1(n10076), .A2(n9693), .ZN(n6938) );
  NAND2_X2 U6854 ( .A1(n10075), .A2(n10082), .ZN(n6939) );
  NAND2_X2 U6855 ( .A1(n6938), .A2(n6939), .ZN(n10077) );
  OR2_X4 U6856 ( .A1(n10077), .A2(n10085), .ZN(n12399) );
  AOI21_X2 U6857 ( .B1(n10025), .B2(n10024), .A(n10023), .ZN(n10042) );
  OAI22_X1 U6858 ( .A1(n6970), .A2(n7108), .B1(n9819), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[17]) );
  NOR2_X1 U6859 ( .A1(pipeline_rs1_data_bypassed[19]), .A2(n9463), .ZN(n10959)
         );
  INV_X4 U6860 ( .A(pipeline_rs1_data_bypassed[17]), .ZN(n12470) );
  AND2_X2 U6861 ( .A1(n8086), .A2(n8087), .ZN(n8085) );
  AND2_X2 U6862 ( .A1(n8888), .A2(n8889), .ZN(n8887) );
  INV_X1 U6863 ( .A(n9667), .ZN(n12994) );
  OAI22_X1 U6864 ( .A1(n6604), .A2(n12565), .B1(n12064), .B2(n12273), .ZN(
        n11799) );
  AOI221_X1 U6865 ( .B1(n9471), .B2(n6610), .C1(n12276), .C2(n6604), .A(n11368), .ZN(n11946) );
  INV_X2 U6866 ( .A(n9834), .ZN(n9831) );
  OAI221_X1 U6867 ( .B1(n7006), .B2(n11405), .C1(n6997), .C2(n11404), .A(
        n11396), .ZN(n11679) );
  NAND2_X1 U6868 ( .A1(n6618), .A2(n11405), .ZN(n11574) );
  OAI22_X1 U6869 ( .A1(n9447), .A2(n7126), .B1(n12862), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[26]) );
  OAI22_X1 U6870 ( .A1(n9447), .A2(n7125), .B1(n12860), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[27]) );
  NOR2_X1 U6871 ( .A1(n12509), .A2(n9486), .ZN(n12510) );
  AND4_X2 U6872 ( .A1(n9263), .A2(n9264), .A3(n9265), .A4(n9266), .ZN(n7101)
         );
  AND3_X2 U6873 ( .A1(n6992), .A2(n6991), .A3(n6990), .ZN(n9266) );
  NAND2_X1 U6874 ( .A1(pipeline_regfile_data[415]), .A2(n9331), .ZN(n9277) );
  NAND2_X2 U6875 ( .A1(n9388), .A2(n9891), .ZN(n9883) );
  OAI22_X2 U6876 ( .A1(n734), .A2(n9445), .B1(n12462), .B2(n9443), .ZN(
        pipeline_alu_src_a[19]) );
  INV_X1 U6877 ( .A(n9888), .ZN(n9889) );
  AOI221_X1 U6878 ( .B1(pipeline_regfile_data[105]), .B2(n8248), .C1(
        pipeline_regfile_data[41]), .C2(n8253), .A(n7522), .ZN(n7521) );
  AOI221_X1 U6879 ( .B1(pipeline_regfile_data[107]), .B2(n8248), .C1(
        pipeline_regfile_data[43]), .C2(n8253), .A(n7586), .ZN(n7585) );
  AND4_X2 U6880 ( .A1(n7952), .A2(n7953), .A3(n7954), .A4(n7955), .ZN(n7123)
         );
  AOI221_X1 U6881 ( .B1(pipeline_regfile_data[118]), .B2(n8246), .C1(
        pipeline_regfile_data[54]), .C2(n8252), .A(n7937), .ZN(n7936) );
  INV_X2 U6882 ( .A(n8431), .ZN(n8430) );
  NAND2_X2 U6883 ( .A1(n9904), .A2(n9903), .ZN(n9895) );
  AOI221_X1 U6884 ( .B1(n12172), .B2(n11376), .C1(n11375), .C2(
        pipeline_alu_src_b[16]), .A(n11374), .ZN(n11381) );
  NOR2_X1 U6885 ( .A1(pipeline_alu_src_b[16]), .A2(n12357), .ZN(n11371) );
  OAI221_X1 U6886 ( .B1(n7214), .B2(n10302), .C1(n12413), .C2(n9467), .A(
        n10301), .ZN(n10422) );
  NOR2_X1 U6887 ( .A1(n12413), .A2(n9484), .ZN(n12414) );
  INV_X2 U6888 ( .A(n12399), .ZN(n10078) );
  INV_X2 U6889 ( .A(n8425), .ZN(n8424) );
  INV_X4 U6890 ( .A(n9322), .ZN(n9324) );
  INV_X4 U6891 ( .A(pipeline_rs1_data_bypassed[31]), .ZN(n12413) );
  NAND2_X2 U6892 ( .A1(n6369), .A2(n9395), .ZN(n6944) );
  OR2_X1 U6893 ( .A1(n9487), .A2(n12457), .ZN(n6945) );
  OR2_X1 U6894 ( .A1(n1504), .A2(n6661), .ZN(n6946) );
  NAND3_X2 U6895 ( .A1(n6945), .A2(n6946), .A3(n12456), .ZN(
        pipeline_PCmux_base[21]) );
  OAI221_X2 U6896 ( .B1(n9488), .B2(n12445), .C1(n1507), .C2(n6661), .A(n12444), .ZN(pipeline_PCmux_base[24]) );
  AOI221_X1 U6897 ( .B1(pipeline_md_N65), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[2]), .A(n12744), .ZN(n12745) );
  NAND2_X1 U6898 ( .A1(n11695), .A2(pipeline_alu_src_b[21]), .ZN(n11696) );
  NOR2_X1 U6899 ( .A1(pipeline_alu_src_b[21]), .A2(n12357), .ZN(n11678) );
  INV_X2 U6900 ( .A(pipeline_alu_src_b[21]), .ZN(n9816) );
  AND4_X2 U6901 ( .A1(n7888), .A2(n7889), .A3(n7890), .A4(n7891), .ZN(n7129)
         );
  AOI221_X1 U6902 ( .B1(pipeline_regfile_data[117]), .B2(n8246), .C1(
        pipeline_regfile_data[53]), .C2(n8252), .A(n7905), .ZN(n7904) );
  AOI221_X1 U6903 ( .B1(pipeline_regfile_data[121]), .B2(n8246), .C1(
        pipeline_regfile_data[57]), .C2(n8252), .A(n8033), .ZN(n8032) );
  INV_X4 U6904 ( .A(n12411), .ZN(n12408) );
  INV_X2 U6905 ( .A(n9267), .ZN(n6992) );
  NOR3_X4 U6906 ( .A1(n6786), .A2(n9585), .A3(n9584), .ZN(n9588) );
  INV_X4 U6907 ( .A(n7987), .ZN(n7030) );
  AND2_X2 U6908 ( .A1(n7257), .A2(n7258), .ZN(n7256) );
  NAND2_X1 U6909 ( .A1(pipeline_regfile_data[490]), .A2(n8254), .ZN(n7548) );
  NAND2_X1 U6910 ( .A1(pipeline_regfile_data[487]), .A2(n8254), .ZN(n7452) );
  AND2_X1 U6911 ( .A1(pipeline_PC_DX[12]), .A2(n9336), .ZN(n6947) );
  AND2_X1 U6912 ( .A1(pipeline_handler_PC[12]), .A2(n6630), .ZN(n6948) );
  NOR3_X2 U6913 ( .A1(n6947), .A2(n6948), .A3(n12490), .ZN(n12491) );
  OR2_X1 U6914 ( .A1(n9487), .A2(n12492), .ZN(n6949) );
  OR2_X1 U6915 ( .A1(n1495), .A2(n6661), .ZN(n6950) );
  NAND3_X2 U6916 ( .A1(n6949), .A2(n6950), .A3(n12491), .ZN(
        pipeline_PCmux_base[12]) );
  OAI21_X4 U6917 ( .B1(n9588), .B2(n9587), .A(n9586), .ZN(n12599) );
  NOR2_X1 U6918 ( .A1(n12489), .A2(n9485), .ZN(n12490) );
  NOR2_X2 U6919 ( .A1(n6951), .A2(n6952), .ZN(n9880) );
  AND2_X1 U6920 ( .A1(n9867), .A2(n9869), .ZN(n6951) );
  NAND2_X2 U6921 ( .A1(n9394), .A2(n6778), .ZN(n6952) );
  INV_X2 U6922 ( .A(n9882), .ZN(n9875) );
  OAI22_X1 U6923 ( .A1(n12967), .A2(n10055), .B1(n9447), .B2(n7148), .ZN(n6987) );
  AOI221_X1 U6924 ( .B1(n11882), .B2(n6611), .C1(n12062), .C2(n11881), .A(
        n11880), .ZN(n11889) );
  NAND2_X1 U6925 ( .A1(n12276), .A2(n6612), .ZN(n11718) );
  NAND2_X1 U6926 ( .A1(n9489), .A2(n6611), .ZN(n11870) );
  NAND2_X2 U6927 ( .A1(n12561), .A2(n12557), .ZN(n12542) );
  OAI22_X2 U6928 ( .A1(n8214), .A2(n12562), .B1(n598), .B2(n12561), .ZN(
        pipeline_PCmux_offset[4]) );
  NAND3_X2 U6929 ( .A1(n6791), .A2(n9898), .A3(n9897), .ZN(n9908) );
  AND4_X2 U6930 ( .A1(n8175), .A2(n8176), .A3(n8177), .A4(n8178), .ZN(n7137)
         );
  AOI221_X1 U6931 ( .B1(n11729), .B2(n6620), .C1(n12062), .C2(n11728), .A(
        n11727), .ZN(n11736) );
  NAND2_X1 U6932 ( .A1(n12276), .A2(n6621), .ZN(n12131) );
  NAND2_X1 U6933 ( .A1(n9489), .A2(n6621), .ZN(n11716) );
  AND2_X2 U6934 ( .A1(n7608), .A2(n7609), .ZN(n7607) );
  INV_X2 U6935 ( .A(n9933), .ZN(n9935) );
  OAI22_X2 U6936 ( .A1(n11656), .A2(n9453), .B1(n6924), .B2(n9450), .ZN(n9933)
         );
  AOI221_X1 U6937 ( .B1(n12268), .B2(n12363), .C1(n12267), .C2(
        pipeline_alu_src_a[2]), .A(n12266), .ZN(n12287) );
  NOR2_X1 U6938 ( .A1(pipeline_alu_src_a[2]), .A2(n12357), .ZN(n12263) );
  NAND2_X1 U6939 ( .A1(n11869), .A2(pipeline_alu_src_a[2]), .ZN(n11400) );
  NAND2_X1 U6940 ( .A1(n9471), .A2(pipeline_alu_src_a[2]), .ZN(n12369) );
  NOR2_X1 U6941 ( .A1(pipeline_alu_src_a[2]), .A2(n12565), .ZN(n11166) );
  OAI21_X2 U6942 ( .B1(n9909), .B2(n9908), .A(n9907), .ZN(n9921) );
  OAI221_X1 U6943 ( .B1(n11474), .B2(n11373), .C1(n11372), .C2(n11407), .A(
        n12659), .ZN(n11374) );
  AOI221_X1 U6944 ( .B1(n9471), .B2(n11546), .C1(n12276), .C2(n11474), .A(
        n11473), .ZN(n12647) );
  AOI221_X1 U6945 ( .B1(n9471), .B2(n11474), .C1(n12276), .C2(n11414), .A(
        n11413), .ZN(n12014) );
  OAI221_X1 U6946 ( .B1(n11414), .B2(n11574), .C1(n11474), .C2(n11572), .A(
        n11156), .ZN(n12281) );
  OAI221_X1 U6947 ( .B1(n11474), .B2(n11574), .C1(n11546), .C2(n11572), .A(
        n11332), .ZN(n11877) );
  OAI22_X1 U6948 ( .A1(n11573), .A2(n12565), .B1(n11474), .B2(n9401), .ZN(
        n11436) );
  INV_X1 U6949 ( .A(n9836), .ZN(n9838) );
  INV_X4 U6950 ( .A(pipeline_alu_src_a[16]), .ZN(n11474) );
  INV_X4 U6951 ( .A(pipeline_rs1_data_bypassed[4]), .ZN(n12522) );
  INV_X4 U6952 ( .A(n13161), .ZN(n6953) );
  AOI221_X1 U6953 ( .B1(pipeline_md_N29), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[0]), .A(n10267), .ZN(n10268) );
  AOI221_X1 U6954 ( .B1(n9483), .B2(pipeline_rs1_data_bypassed[0]), .C1(
        pipeline_PC_DX[0]), .C2(n6969), .A(n12540), .ZN(n12541) );
  NAND2_X1 U6955 ( .A1(n11869), .A2(pipeline_alu_src_a[0]), .ZN(n11341) );
  OAI221_X1 U6956 ( .B1(n6632), .B2(n11404), .C1(pipeline_alu_src_a[0]), .C2(
        n11405), .A(n11167), .ZN(n11507) );
  NAND2_X1 U6957 ( .A1(n9489), .A2(pipeline_alu_src_a[0]), .ZN(n11610) );
  MUX2_X1 U6958 ( .A(pipeline_alu_src_a[0]), .B(n6632), .S(n11404), .Z(n11406)
         );
  OAI221_X1 U6959 ( .B1(n594), .B2(n12561), .C1(n693), .C2(n12557), .A(n12553), 
        .ZN(pipeline_PCmux_offset[11]) );
  NOR2_X2 U6960 ( .A1(n12492), .A2(n9494), .ZN(n6954) );
  NOR2_X2 U6961 ( .A1(n9493), .A2(n9354), .ZN(n6955) );
  OR2_X2 U6962 ( .A1(n6954), .A2(n6955), .ZN(n5959) );
  INV_X8 U6963 ( .A(n9378), .ZN(imem_haddr[27]) );
  AOI221_X1 U6964 ( .B1(pipeline_md_N68), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[5]), .A(n12738), .ZN(n12739) );
  OAI221_X1 U6965 ( .B1(n11280), .B2(n636), .C1(n11279), .C2(n9467), .A(n11278), .ZN(n12622) );
  NAND2_X2 U6966 ( .A1(n12561), .A2(n12557), .ZN(n6958) );
  OR2_X4 U6967 ( .A1(n7056), .A2(n7057), .ZN(pipeline_rs1_data_bypassed[3]) );
  NOR2_X2 U6968 ( .A1(n12967), .A2(n9784), .ZN(n7057) );
  INV_X1 U6969 ( .A(ext_interrupts[7]), .ZN(n6959) );
  INV_X1 U6970 ( .A(n6959), .ZN(n6960) );
  OAI221_X1 U6971 ( .B1(n7185), .B2(n10689), .C1(n12509), .C2(n9467), .A(n4130), .ZN(n11892) );
  INV_X4 U6972 ( .A(n6987), .ZN(n9707) );
  INV_X4 U6973 ( .A(n9385), .ZN(n9891) );
  AOI22_X2 U6974 ( .A1(n6600), .A2(n9457), .B1(pipeline_alu_src_a[4]), .B2(
        n9452), .ZN(n9385) );
  AND2_X2 U6975 ( .A1(pipeline_PC_DX[14]), .A2(n9336), .ZN(n6961) );
  AND2_X1 U6976 ( .A1(pipeline_handler_PC[14]), .A2(n6630), .ZN(n6962) );
  NOR3_X1 U6977 ( .A1(n6961), .A2(n6962), .A3(n12482), .ZN(n12483) );
  OR2_X1 U6978 ( .A1(n9488), .A2(n12484), .ZN(n6963) );
  OR2_X1 U6979 ( .A1(n1497), .A2(n6661), .ZN(n6964) );
  NAND3_X2 U6980 ( .A1(n6963), .A2(n6964), .A3(n12483), .ZN(
        pipeline_PCmux_base[14]) );
  NOR2_X1 U6981 ( .A1(n12481), .A2(n9485), .ZN(n12482) );
  AOI221_X1 U6982 ( .B1(n11584), .B2(n11583), .C1(n11582), .C2(n6614), .A(
        n11581), .ZN(n11592) );
  NAND2_X1 U6983 ( .A1(n12276), .A2(n6614), .ZN(n11722) );
  NAND2_X1 U6984 ( .A1(n9489), .A2(n6614), .ZN(n11569) );
  OAI22_X1 U6985 ( .A1(pipeline_alu_src_a[14]), .A2(n12565), .B1(n6614), .B2(
        n9401), .ZN(n11168) );
  NAND2_X1 U6986 ( .A1(pipeline_PC_DX[16]), .A2(n9336), .ZN(n6965) );
  NAND2_X1 U6987 ( .A1(pipeline_handler_PC[16]), .A2(n6630), .ZN(n6966) );
  AND3_X2 U6988 ( .A1(n6965), .A2(n6966), .A3(n6577), .ZN(n12475) );
  OR2_X1 U6989 ( .A1(n9488), .A2(n12476), .ZN(n6967) );
  OR2_X1 U6990 ( .A1(n1499), .A2(n6661), .ZN(n6968) );
  INV_X16 U6991 ( .A(n9483), .ZN(n9485) );
  AOI221_X1 U6992 ( .B1(pipeline_md_N56), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[27]), .A(n10453), .ZN(n10454) );
  NOR2_X1 U6993 ( .A1(pipeline_rs1_data_bypassed[27]), .A2(n9463), .ZN(n10476)
         );
  NAND2_X1 U6994 ( .A1(n9471), .A2(n6602), .ZN(n12212) );
  NAND2_X1 U6995 ( .A1(n12276), .A2(n6603), .ZN(n12308) );
  NAND2_X1 U6996 ( .A1(n9489), .A2(n6602), .ZN(n12175) );
  NAND2_X1 U6997 ( .A1(n11869), .A2(n6602), .ZN(n12651) );
  OAI221_X1 U6998 ( .B1(n7213), .B2(n10633), .C1(n12505), .C2(n9467), .A(n3718), .ZN(n11999) );
  NOR2_X1 U6999 ( .A1(n12505), .A2(n9485), .ZN(n12506) );
  INV_X8 U7000 ( .A(n10798), .ZN(imem_haddr[26]) );
  INV_X8 U7001 ( .A(n10451), .ZN(imem_haddr[28]) );
  INV_X8 U7002 ( .A(n10387), .ZN(imem_haddr[29]) );
  INV_X8 U7003 ( .A(n6953), .ZN(imem_haddr[30]) );
  INV_X8 U7004 ( .A(n12563), .ZN(imem_haddr[31]) );
  NOR2_X2 U7005 ( .A1(n12442), .A2(n9484), .ZN(n12443) );
  NAND2_X1 U7006 ( .A1(n12552), .A2(n12551), .ZN(pipeline_PCmux_offset[12]) );
  NAND2_X1 U7007 ( .A1(n12552), .A2(n12547), .ZN(pipeline_PCmux_offset[17]) );
  NAND2_X1 U7008 ( .A1(n9391), .A2(n10258), .ZN(n6970) );
  INV_X4 U7009 ( .A(n6942), .ZN(n9439) );
  INV_X4 U7010 ( .A(n6942), .ZN(n9440) );
  NAND2_X1 U7011 ( .A1(n12552), .A2(n12548), .ZN(pipeline_PCmux_offset[14]) );
  NAND2_X1 U7012 ( .A1(n12552), .A2(n12549), .ZN(pipeline_PCmux_offset[13]) );
  NOR2_X2 U7013 ( .A1(n12530), .A2(n9486), .ZN(n12531) );
  INV_X4 U7014 ( .A(pipeline_alu_src_a[9]), .ZN(n6971) );
  INV_X4 U7015 ( .A(n6971), .ZN(n6972) );
  INV_X1 U7016 ( .A(n6971), .ZN(n6973) );
  INV_X1 U7017 ( .A(n9388), .ZN(n9892) );
  INV_X4 U7018 ( .A(pipeline_alu_src_b[1]), .ZN(n6974) );
  INV_X4 U7019 ( .A(n6974), .ZN(n6975) );
  INV_X1 U7020 ( .A(n6974), .ZN(n6976) );
  NAND2_X2 U7021 ( .A1(n9724), .A2(n9723), .ZN(n9392) );
  AOI21_X2 U7022 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9863) );
  INV_X4 U7023 ( .A(n9333), .ZN(n9329) );
  INV_X1 U7024 ( .A(n9333), .ZN(n9332) );
  INV_X1 U7025 ( .A(n9333), .ZN(n9331) );
  AOI221_X1 U7026 ( .B1(pipeline_dmem_type_2_), .B2(n601), .C1(n6784), .C2(
        n713), .A(dmem_hsize[1]), .ZN(n9680) );
  NOR2_X2 U7027 ( .A1(n12500), .A2(n9494), .ZN(n6977) );
  NOR2_X2 U7028 ( .A1(n9493), .A2(n9358), .ZN(n6978) );
  OR2_X2 U7029 ( .A1(n6977), .A2(n6978), .ZN(n5961) );
  OAI22_X1 U7030 ( .A1(n6970), .A2(n7109), .B1(n9997), .B2(n9441), .ZN(n6979)
         );
  AND4_X4 U7031 ( .A1(n9007), .A2(n9008), .A3(n9009), .A4(n9010), .ZN(n7109)
         );
  OAI22_X1 U7032 ( .A1(n738), .A2(n9445), .B1(n12446), .B2(n9443), .ZN(n6980)
         );
  AND2_X1 U7033 ( .A1(pipeline_regfile_data[932]), .A2(n6767), .ZN(n6981) );
  AND2_X1 U7034 ( .A1(pipeline_regfile_data[676]), .A2(n6764), .ZN(n6982) );
  NOR3_X2 U7035 ( .A1(n6981), .A2(n6982), .A3(n8405), .ZN(n8404) );
  OR2_X4 U7036 ( .A1(n8406), .A2(n9305), .ZN(n6983) );
  OR2_X4 U7037 ( .A1(n8407), .A2(n9306), .ZN(n6984) );
  NAND2_X2 U7038 ( .A1(n6983), .A2(n6984), .ZN(n8405) );
  AND2_X4 U7039 ( .A1(n8416), .A2(n8417), .ZN(n8406) );
  AND2_X2 U7040 ( .A1(n8408), .A2(n8409), .ZN(n8407) );
  AND2_X4 U7041 ( .A1(pipeline_PC_DX[6]), .A2(n6969), .ZN(n6985) );
  AND2_X1 U7042 ( .A1(pipeline_handler_PC[6]), .A2(n6630), .ZN(n6986) );
  NOR3_X2 U7043 ( .A1(n6985), .A2(n6986), .A3(n12514), .ZN(n12515) );
  NOR2_X1 U7044 ( .A1(n12513), .A2(n9486), .ZN(n12514) );
  OAI22_X2 U7045 ( .A1(n12967), .A2(n6638), .B1(n9447), .B2(n7148), .ZN(
        pipeline_rs2_data_bypassed[3]) );
  AND2_X1 U7046 ( .A1(pipeline_regfile_data[931]), .A2(n6767), .ZN(n6988) );
  AND2_X1 U7047 ( .A1(pipeline_regfile_data[675]), .A2(n6764), .ZN(n6989) );
  NOR3_X2 U7048 ( .A1(n6988), .A2(n6989), .A3(n8376), .ZN(n8375) );
  NAND2_X1 U7049 ( .A1(pipeline_regfile_data[959]), .A2(n6767), .ZN(n6990) );
  NAND2_X1 U7050 ( .A1(pipeline_regfile_data[703]), .A2(n6764), .ZN(n6991) );
  AND2_X1 U7051 ( .A1(pipeline_regfile_data[929]), .A2(n6767), .ZN(n6993) );
  AND2_X1 U7052 ( .A1(pipeline_regfile_data[673]), .A2(n6764), .ZN(n6994) );
  OR2_X4 U7053 ( .A1(n732), .A2(n9445), .ZN(n6995) );
  OR2_X4 U7054 ( .A1(n12470), .A2(n9443), .ZN(n6996) );
  NAND2_X1 U7055 ( .A1(n11869), .A2(pipeline_alu_src_a[17]), .ZN(n11618) );
  OAI22_X1 U7056 ( .A1(pipeline_alu_src_a[17]), .A2(n12565), .B1(
        pipeline_alu_src_a[14]), .B2(n9400), .ZN(n11413) );
  NAND2_X1 U7057 ( .A1(n9471), .A2(pipeline_alu_src_a[17]), .ZN(n9748) );
  NAND2_X1 U7058 ( .A1(n9489), .A2(pipeline_alu_src_a[17]), .ZN(n11397) );
  INV_X4 U7059 ( .A(n12635), .ZN(n6997) );
  INV_X1 U7060 ( .A(pipeline_alu_src_a[30]), .ZN(n12635) );
  OAI22_X2 U7061 ( .A1(n745), .A2(n9445), .B1(n12418), .B2(n9443), .ZN(
        pipeline_alu_src_a[30]) );
  AND2_X2 U7062 ( .A1(pipeline_regfile_N12), .A2(pipeline_regfile_N13), .ZN(
        n7170) );
  AOI221_X1 U7063 ( .B1(n603), .B2(pipeline_rs1_data_bypassed[0]), .C1(
        pipeline_regfile_N12), .C2(pipeline_dmem_type_2_), .A(n11276), .ZN(
        n11277) );
  XNOR2_X1 U7064 ( .A(n12990), .B(pipeline_regfile_N12), .ZN(n9645) );
  OAI22_X1 U7065 ( .A1(n9439), .A2(n7070), .B1(n12962), .B2(n9393), .ZN(n6998)
         );
  OAI22_X2 U7066 ( .A1(n9440), .A2(n7070), .B1(n12962), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[4]) );
  NAND2_X1 U7067 ( .A1(pipeline_regfile_data[945]), .A2(n6728), .ZN(n6999) );
  INV_X4 U7068 ( .A(n7764), .ZN(n7001) );
  NAND2_X1 U7069 ( .A1(pipeline_regfile_N18), .A2(pipeline_regfile_N19), .ZN(
        n7002) );
  INV_X2 U7070 ( .A(n7002), .ZN(n7003) );
  OAI22_X1 U7071 ( .A1(n12962), .A2(n10055), .B1(n7061), .B2(n7071), .ZN(n7004) );
  OAI22_X2 U7072 ( .A1(n12962), .A2(n10055), .B1(n9447), .B2(n7071), .ZN(
        pipeline_rs2_data_bypassed[4]) );
  INV_X1 U7073 ( .A(n6744), .ZN(n9452) );
  OAI22_X1 U7074 ( .A1(n746), .A2(n9786), .B1(n12413), .B2(n9443), .ZN(n7005)
         );
  OAI22_X1 U7075 ( .A1(n746), .A2(n9786), .B1(n12413), .B2(n9443), .ZN(n7006)
         );
  NOR2_X1 U7076 ( .A1(pipeline_alu_src_b[20]), .A2(n12357), .ZN(n11611) );
  AND4_X2 U7077 ( .A1(n7633), .A2(n7634), .A3(n7635), .A4(n7636), .ZN(n7118)
         );
  NAND2_X1 U7078 ( .A1(pipeline_inst_DX[10]), .A2(n9712), .ZN(n7007) );
  NAND2_X2 U7079 ( .A1(pipeline_rs2_data_bypassed[3]), .A2(n9449), .ZN(n7008)
         );
  NAND2_X1 U7080 ( .A1(n9398), .A2(n7009), .ZN(n12774) );
  NAND2_X1 U7081 ( .A1(n7084), .A2(n7009), .ZN(n11372) );
  OAI221_X1 U7082 ( .B1(n9509), .B2(n11876), .C1(n7009), .C2(n11583), .A(
        n11530), .ZN(n12127) );
  OAI221_X1 U7083 ( .B1(n7009), .B2(n12362), .C1(n9399), .C2(n12013), .A(
        n12012), .ZN(n12068) );
  NAND2_X1 U7084 ( .A1(n11953), .A2(n7009), .ZN(n11986) );
  NAND2_X1 U7085 ( .A1(n11756), .A2(n7009), .ZN(n11810) );
  NAND2_X1 U7086 ( .A1(n12165), .A2(n7009), .ZN(n12168) );
  NAND2_X1 U7087 ( .A1(n11828), .A2(n7009), .ZN(n11886) );
  NAND2_X1 U7088 ( .A1(n7009), .A2(n9399), .ZN(n12776) );
  OAI221_X1 U7089 ( .B1(n11653), .B2(n9509), .C1(n7009), .C2(n11652), .A(
        n11651), .ZN(n12218) );
  OAI221_X1 U7090 ( .B1(n7009), .B2(n12268), .C1(n9399), .C2(n11755), .A(
        n11509), .ZN(n12085) );
  OAI221_X1 U7091 ( .B1(n7009), .B2(n12126), .C1(n9399), .C2(n11827), .A(
        n11586), .ZN(n12160) );
  OAI221_X1 U7092 ( .B1(n11946), .B2(n9509), .C1(n7009), .C2(n7084), .A(n11945), .ZN(n11993) );
  NAND2_X1 U7093 ( .A1(n12174), .A2(n7009), .ZN(n11613) );
  NAND2_X1 U7094 ( .A1(n11674), .A2(n7009), .ZN(n11733) );
  INV_X1 U7095 ( .A(n10009), .ZN(n9810) );
  AOI211_X2 U7096 ( .C1(n9863), .C2(n9900), .A(n9862), .B(n9861), .ZN(n9922)
         );
  AOI21_X2 U7097 ( .B1(n9610), .B2(n9609), .A(n12148), .ZN(n9611) );
  AOI221_X1 U7098 ( .B1(pipeline_regfile_data[706]), .B2(n6734), .C1(
        pipeline_regfile_data[898]), .C2(n6733), .A(n7307), .ZN(n7282) );
  AND4_X4 U7099 ( .A1(n8016), .A2(n8017), .A3(n8018), .A4(n8019), .ZN(n7124)
         );
  AND4_X4 U7100 ( .A1(n7792), .A2(n7793), .A3(n7794), .A4(n7795), .ZN(n7132)
         );
  AND4_X4 U7101 ( .A1(n7824), .A2(n7825), .A3(n7826), .A4(n7827), .ZN(n7134)
         );
  AND4_X4 U7102 ( .A1(n7920), .A2(n7921), .A3(n7922), .A4(n7923), .ZN(n7133)
         );
  AOI221_X1 U7103 ( .B1(pipeline_regfile_data[734]), .B2(n6734), .C1(
        pipeline_regfile_data[926]), .C2(n6733), .A(n8201), .ZN(n8176) );
  AND4_X4 U7104 ( .A1(n8849), .A2(n8850), .A3(n8851), .A4(n8852), .ZN(n7106)
         );
  AOI221_X1 U7105 ( .B1(pipeline_regfile_data[718]), .B2(n6773), .C1(
        pipeline_regfile_data[910]), .C2(n6772), .A(n8747), .ZN(n8722) );
  AND4_X4 U7106 ( .A1(n8721), .A2(n8722), .A3(n8723), .A4(n8724), .ZN(n7092)
         );
  AOI221_X1 U7107 ( .B1(n12790), .B2(n12789), .C1(n12788), .C2(n6927), .A(
        n12787), .ZN(n12803) );
  NAND2_X1 U7108 ( .A1(n9471), .A2(pipeline_alu_src_a[4]), .ZN(n12132) );
  NAND2_X1 U7109 ( .A1(n11869), .A2(n6928), .ZN(n12367) );
  AOI221_X1 U7110 ( .B1(n9471), .B2(n6634), .C1(n12276), .C2(n6927), .A(n12275), .ZN(n12277) );
  OAI22_X1 U7111 ( .A1(pipeline_alu_src_a[4]), .A2(n12565), .B1(n6632), .B2(
        n9400), .ZN(n11365) );
  INV_X1 U7112 ( .A(n6928), .ZN(n12792) );
  INV_X4 U7113 ( .A(n8244), .ZN(n8249) );
  INV_X2 U7114 ( .A(n8244), .ZN(n8248) );
  INV_X2 U7115 ( .A(n7015), .ZN(n8264) );
  INV_X2 U7116 ( .A(n6642), .ZN(n8259) );
  INV_X2 U7117 ( .A(n6642), .ZN(n8260) );
  OAI22_X1 U7118 ( .A1(n7082), .A2(n9507), .B1(n12133), .B2(n12582), .ZN(
        n12134) );
  OAI221_X1 U7119 ( .B1(n12582), .B2(n11466), .C1(n9507), .C2(n12087), .A(
        n11465), .ZN(n11470) );
  OAI221_X1 U7120 ( .B1(n12582), .B2(n12017), .C1(n12016), .C2(n9507), .A(
        n12015), .ZN(n12023) );
  OAI221_X1 U7121 ( .B1(n11443), .B2(n12582), .C1(n9507), .C2(n12017), .A(
        n11402), .ZN(n11410) );
  OAI221_X1 U7122 ( .B1(n11532), .B2(n12582), .C1(n12774), .C2(n12164), .A(
        n11531), .ZN(n11538) );
  OAI221_X1 U7123 ( .B1(n12582), .B2(n11944), .C1(n9507), .C2(n11950), .A(
        n11369), .ZN(n11376) );
  AND2_X4 U7124 ( .A1(n9658), .A2(n693), .ZN(n7078) );
  INV_X1 U7125 ( .A(n10388), .ZN(n10098) );
  INV_X2 U7126 ( .A(n9298), .ZN(n9311) );
  AOI221_X2 U7127 ( .B1(pipeline_inst_DX[9]), .B2(n9712), .C1(n9449), .C2(
        pipeline_rs2_data_bypassed[2]), .A(n9711), .ZN(n12265) );
  AOI221_X2 U7128 ( .B1(pipeline_regfile_data[704]), .B2(n6734), .C1(
        pipeline_regfile_data[896]), .C2(n6733), .A(n7244), .ZN(n7218) );
  INV_X4 U7129 ( .A(n8311), .ZN(n7019) );
  NOR4_X2 U7130 ( .A1(n7017), .A2(n7018), .A3(n7019), .A4(n6782), .ZN(n7097)
         );
  AND4_X4 U7131 ( .A1(n9071), .A2(n9072), .A3(n9073), .A4(n9074), .ZN(n7105)
         );
  NOR4_X2 U7132 ( .A1(n7024), .A2(n7025), .A3(n7026), .A4(n6783), .ZN(n7126)
         );
  INV_X4 U7133 ( .A(n8343), .ZN(n7041) );
  INV_X4 U7134 ( .A(n8342), .ZN(n7040) );
  NOR4_X2 U7135 ( .A1(n7038), .A2(n7039), .A3(n7040), .A4(n7041), .ZN(n7138)
         );
  INV_X4 U7136 ( .A(n8468), .ZN(n7045) );
  INV_X4 U7137 ( .A(n8467), .ZN(n7044) );
  NOR4_X2 U7138 ( .A1(n7042), .A2(n7043), .A3(n7044), .A4(n7045), .ZN(n7141)
         );
  AND2_X4 U7139 ( .A1(pipeline_regfile_N16), .A2(pipeline_regfile_N15), .ZN(
        n7164) );
  OAI22_X1 U7140 ( .A1(n6639), .A2(n12824), .B1(n6628), .B2(n12823), .ZN(n6284) );
  NOR2_X2 U7141 ( .A1(n6970), .A2(n6790), .ZN(n7056) );
  INV_X1 U7142 ( .A(n6573), .ZN(n9457) );
  INV_X1 U7143 ( .A(n6573), .ZN(n9459) );
  INV_X2 U7144 ( .A(n6642), .ZN(n8258) );
  INV_X4 U7145 ( .A(n9354), .ZN(imem_haddr[12]) );
  INV_X4 U7146 ( .A(n9358), .ZN(imem_haddr[10]) );
  INV_X4 U7147 ( .A(n9348), .ZN(imem_haddr[15]) );
  INV_X4 U7148 ( .A(n9342), .ZN(imem_haddr[8]) );
  OAI221_X1 U7149 ( .B1(n12099), .B2(n12090), .C1(n6806), .C2(n12089), .A(
        n12659), .ZN(n12091) );
  OAI221_X1 U7150 ( .B1(n12582), .B2(n12164), .C1(n12163), .C2(n9507), .A(
        n12162), .ZN(n12171) );
  INV_X2 U7151 ( .A(n9312), .ZN(n9314) );
  NAND2_X2 U7152 ( .A1(pipeline_alu_N284), .A2(n6812), .ZN(n7059) );
  INV_X4 U7154 ( .A(n8250), .ZN(n8251) );
  INV_X4 U7155 ( .A(n11264), .ZN(n13108) );
  OAI221_X1 U7156 ( .B1(n12582), .B2(n11650), .C1(n12774), .C2(n12221), .A(
        n11609), .ZN(n11615) );
  OAI221_X1 U7157 ( .B1(n11677), .B2(n12582), .C1(n12774), .C2(n12317), .A(
        n11676), .ZN(n11684) );
  OAI221_X1 U7158 ( .B1(n12582), .B2(n11761), .C1(n12774), .C2(n11760), .A(
        n11759), .ZN(n11767) );
  OAI221_X1 U7159 ( .B1(n11832), .B2(n12582), .C1(n9507), .C2(n12581), .A(
        n11831), .ZN(n11839) );
  OAI221_X1 U7160 ( .B1(n12582), .B2(n11950), .C1(n11949), .C2(n9507), .A(
        n11948), .ZN(n11956) );
  OAI221_X1 U7161 ( .B1(n12582), .B2(n12581), .C1(n6811), .C2(n9507), .A(
        n12580), .ZN(n12583) );
  OAI221_X1 U7162 ( .B1(n12582), .B2(n12221), .C1(n6804), .C2(n9507), .A(
        n12220), .ZN(n12222) );
  OAI221_X1 U7163 ( .B1(n12582), .B2(n12317), .C1(n6805), .C2(n9507), .A(
        n12316), .ZN(n12318) );
  OAI221_X1 U7164 ( .B1(n12582), .B2(n12087), .C1(n6800), .C2(n9507), .A(
        n12086), .ZN(n12092) );
  INV_X4 U7165 ( .A(n13111), .ZN(n9528) );
  OAI221_X2 U7166 ( .B1(n10131), .B2(n6807), .C1(n7073), .C2(n7074), .A(n6712), 
        .ZN(n7072) );
  INV_X4 U7167 ( .A(n9446), .ZN(n9445) );
  AND3_X4 U7168 ( .A1(n13097), .A2(n13096), .A3(n13095), .ZN(n7090) );
  OAI22_X2 U7169 ( .A1(n12987), .A2(n10055), .B1(n9447), .B2(n6789), .ZN(
        pipeline_rs2_data_bypassed[0]) );
  INV_X4 U7170 ( .A(n8309), .ZN(n7017) );
  INV_X4 U7171 ( .A(n8310), .ZN(n7018) );
  INV_X2 U7172 ( .A(n7604), .ZN(n7023) );
  INV_X2 U7173 ( .A(n7603), .ZN(n7022) );
  INV_X2 U7174 ( .A(n7601), .ZN(n7020) );
  INV_X2 U7175 ( .A(n7602), .ZN(n7021) );
  INV_X2 U7176 ( .A(n8050), .ZN(n7026) );
  INV_X4 U7177 ( .A(n8048), .ZN(n7024) );
  INV_X4 U7178 ( .A(n8049), .ZN(n7025) );
  INV_X4 U7179 ( .A(n8465), .ZN(n7042) );
  INV_X4 U7180 ( .A(n8466), .ZN(n7043) );
  AOI221_X2 U7181 ( .B1(pipeline_PC_DX[24]), .B2(n9337), .C1(
        pipeline_handler_PC[24]), .C2(n6630), .A(n12443), .ZN(n12444) );
  INV_X2 U7182 ( .A(n7253), .ZN(n7049) );
  INV_X2 U7183 ( .A(n7252), .ZN(n7048) );
  INV_X2 U7184 ( .A(n7250), .ZN(n7046) );
  INV_X2 U7185 ( .A(n7251), .ZN(n7047) );
  INV_X4 U7186 ( .A(n8340), .ZN(n7038) );
  INV_X4 U7187 ( .A(n8341), .ZN(n7039) );
  INV_X2 U7188 ( .A(n7986), .ZN(n7029) );
  INV_X2 U7189 ( .A(n7984), .ZN(n7027) );
  INV_X2 U7190 ( .A(n7985), .ZN(n7028) );
  INV_X2 U7191 ( .A(n7859), .ZN(n7034) );
  INV_X2 U7192 ( .A(n7858), .ZN(n7033) );
  INV_X2 U7193 ( .A(n7856), .ZN(n7031) );
  INV_X2 U7194 ( .A(n7857), .ZN(n7032) );
  INV_X2 U7195 ( .A(n7763), .ZN(n7037) );
  INV_X2 U7196 ( .A(n7761), .ZN(n7035) );
  INV_X2 U7197 ( .A(n7762), .ZN(n7036) );
  AND3_X4 U7198 ( .A1(pipeline_regfile_N14), .A2(n636), .A3(n637), .ZN(n7171)
         );
  AND4_X2 U7199 ( .A1(n8689), .A2(n8690), .A3(n8691), .A4(n8692), .ZN(n7103)
         );
  AOI221_X1 U7200 ( .B1(pipeline_regfile_data[525]), .B2(n6709), .C1(
        pipeline_regfile_data[973]), .C2(n6763), .A(n8718), .ZN(n8689) );
  AND4_X4 U7201 ( .A1(n9231), .A2(n9232), .A3(n9233), .A4(n9234), .ZN(n7115)
         );
  AND4_X4 U7202 ( .A1(n9167), .A2(n9168), .A3(n9169), .A4(n9170), .ZN(n7117)
         );
  AND4_X4 U7203 ( .A1(n8111), .A2(n8112), .A3(n8113), .A4(n8114), .ZN(n7136)
         );
  AND4_X4 U7204 ( .A1(n7569), .A2(n7570), .A3(n7571), .A4(n7572), .ZN(n7102)
         );
  AOI221_X1 U7205 ( .B1(pipeline_regfile_data[715]), .B2(n6734), .C1(
        pipeline_regfile_data[907]), .C2(n6733), .A(n7595), .ZN(n7570) );
  AND4_X2 U7206 ( .A1(n8625), .A2(n8626), .A3(n8627), .A4(n8628), .ZN(n7146)
         );
  AND4_X4 U7207 ( .A1(n8207), .A2(n8208), .A3(n8209), .A4(n8210), .ZN(n7143)
         );
  INV_X2 U7208 ( .A(n9143), .ZN(n7150) );
  OAI22_X1 U7209 ( .A1(n6639), .A2(n10108), .B1(n638), .B2(n12823), .ZN(n6280)
         );
  OAI22_X1 U7210 ( .A1(n6639), .A2(n10112), .B1(n636), .B2(n12823), .ZN(n6278)
         );
  OAI22_X1 U7211 ( .A1(n6639), .A2(n10104), .B1(n713), .B2(n12823), .ZN(n6293)
         );
  OAI22_X1 U7212 ( .A1(n6639), .A2(n10115), .B1(n603), .B2(n12823), .ZN(n6277)
         );
  OAI22_X1 U7213 ( .A1(n6639), .A2(n10106), .B1(n595), .B2(n12823), .ZN(n6265)
         );
  OAI22_X1 U7214 ( .A1(n6639), .A2(n10105), .B1(n594), .B2(n12823), .ZN(n6263)
         );
  OAI22_X1 U7215 ( .A1(n6639), .A2(n10107), .B1(n596), .B2(n12823), .ZN(n6267)
         );
  OAI22_X1 U7216 ( .A1(n6639), .A2(n10122), .B1(n10338), .B2(n12823), .ZN(
        n6289) );
  OAI22_X1 U7217 ( .A1(n6639), .A2(n10110), .B1(n9270), .B2(n12823), .ZN(n6282) );
  OAI22_X1 U7218 ( .A1(n6639), .A2(n10109), .B1(n9279), .B2(n12823), .ZN(n6281) );
  OAI22_X1 U7219 ( .A1(n6639), .A2(n10111), .B1(n637), .B2(n12823), .ZN(n6279)
         );
  OAI22_X1 U7220 ( .A1(n6639), .A2(n10117), .B1(n602), .B2(n12823), .ZN(n6275)
         );
  OAI22_X1 U7221 ( .A1(n6639), .A2(n10113), .B1(n598), .B2(n12823), .ZN(n6271)
         );
  OAI22_X1 U7222 ( .A1(n6639), .A2(n10114), .B1(n597), .B2(n12823), .ZN(n6269)
         );
  OAI22_X1 U7223 ( .A1(n6639), .A2(n10121), .B1(n10236), .B2(n12823), .ZN(
        n6290) );
  OAI22_X1 U7224 ( .A1(n1162), .A2(n9530), .B1(n1911), .B2(n6688), .ZN(n6143)
         );
  OAI22_X1 U7225 ( .A1(n1256), .A2(n6689), .B1(n1911), .B2(n6659), .ZN(n6082)
         );
  OAI22_X1 U7226 ( .A1(n1288), .A2(n9529), .B1(n1911), .B2(n6702), .ZN(n6175)
         );
  OAI22_X1 U7227 ( .A1(n1224), .A2(n3683), .B1(n1911), .B2(n6703), .ZN(n6080)
         );
  AND3_X1 U7228 ( .A1(dmem_hsize[0]), .A2(n13096), .A3(n7064), .ZN(n7179) );
  MUX2_X1 U7229 ( .A(pipeline_regfile_data[506]), .B(n9417), .S(n6644), .Z(
        n4767) );
  MUX2_X1 U7230 ( .A(pipeline_regfile_data[474]), .B(n13002), .S(n6645), .Z(
        n4766) );
  MUX2_X1 U7231 ( .A(pipeline_regfile_data[442]), .B(n9417), .S(n6646), .Z(
        n4765) );
  MUX2_X1 U7232 ( .A(pipeline_regfile_data[410]), .B(n13002), .S(n6647), .Z(
        n4764) );
  MUX2_X1 U7233 ( .A(pipeline_regfile_data[378]), .B(n9417), .S(n6648), .Z(
        n4763) );
  MUX2_X1 U7234 ( .A(pipeline_regfile_data[346]), .B(n13002), .S(n6653), .Z(
        n4762) );
  MUX2_X1 U7235 ( .A(pipeline_regfile_data[250]), .B(n9417), .S(n6649), .Z(
        n4759) );
  MUX2_X1 U7236 ( .A(pipeline_regfile_data[218]), .B(n13002), .S(n6650), .Z(
        n4758) );
  MUX2_X1 U7237 ( .A(pipeline_regfile_data[186]), .B(n9417), .S(n6651), .Z(
        n4757) );
  MUX2_X1 U7238 ( .A(pipeline_regfile_data[154]), .B(n13002), .S(n6652), .Z(
        n4756) );
  MUX2_X1 U7239 ( .A(pipeline_regfile_data[122]), .B(n9417), .S(n6654), .Z(
        n4755) );
  MUX2_X1 U7240 ( .A(pipeline_regfile_data[90]), .B(n13002), .S(n6655), .Z(
        n4754) );
  MUX2_X1 U7241 ( .A(pipeline_regfile_data[500]), .B(n13008), .S(n6644), .Z(
        n4953) );
  MUX2_X1 U7242 ( .A(pipeline_regfile_data[468]), .B(n13008), .S(n6645), .Z(
        n4952) );
  MUX2_X1 U7243 ( .A(pipeline_regfile_data[436]), .B(n13008), .S(n6646), .Z(
        n4951) );
  MUX2_X1 U7244 ( .A(pipeline_regfile_data[404]), .B(n13008), .S(n6647), .Z(
        n4950) );
  MUX2_X1 U7245 ( .A(pipeline_regfile_data[244]), .B(n13008), .S(n6649), .Z(
        n4945) );
  MUX2_X1 U7246 ( .A(pipeline_regfile_data[212]), .B(n13008), .S(n6650), .Z(
        n4944) );
  MUX2_X1 U7247 ( .A(pipeline_regfile_data[180]), .B(n13008), .S(n6651), .Z(
        n4943) );
  MUX2_X1 U7248 ( .A(pipeline_regfile_data[148]), .B(n13008), .S(n6652), .Z(
        n4942) );
  MUX2_X1 U7249 ( .A(pipeline_regfile_data[497]), .B(n13011), .S(n6644), .Z(
        n5046) );
  MUX2_X1 U7250 ( .A(pipeline_regfile_data[465]), .B(n13011), .S(n6645), .Z(
        n5045) );
  MUX2_X1 U7251 ( .A(pipeline_regfile_data[433]), .B(n13011), .S(n6646), .Z(
        n5044) );
  MUX2_X1 U7252 ( .A(pipeline_regfile_data[401]), .B(n13011), .S(n6647), .Z(
        n5043) );
  MUX2_X1 U7253 ( .A(pipeline_regfile_data[369]), .B(n13011), .S(n6648), .Z(
        n5042) );
  MUX2_X1 U7254 ( .A(pipeline_regfile_data[241]), .B(n13011), .S(n6649), .Z(
        n5038) );
  MUX2_X1 U7255 ( .A(pipeline_regfile_data[209]), .B(n13011), .S(n6650), .Z(
        n5037) );
  MUX2_X1 U7256 ( .A(pipeline_regfile_data[177]), .B(n13011), .S(n6651), .Z(
        n5036) );
  MUX2_X1 U7257 ( .A(pipeline_regfile_data[145]), .B(n13011), .S(n6652), .Z(
        n5035) );
  MUX2_X1 U7258 ( .A(pipeline_regfile_data[504]), .B(n9419), .S(n6644), .Z(
        n4829) );
  MUX2_X1 U7259 ( .A(pipeline_regfile_data[472]), .B(n13004), .S(n6645), .Z(
        n4828) );
  MUX2_X1 U7260 ( .A(pipeline_regfile_data[440]), .B(n9419), .S(n6646), .Z(
        n4827) );
  MUX2_X1 U7261 ( .A(pipeline_regfile_data[408]), .B(n13004), .S(n6647), .Z(
        n4826) );
  MUX2_X1 U7262 ( .A(pipeline_regfile_data[248]), .B(n9419), .S(n6649), .Z(
        n4821) );
  MUX2_X1 U7263 ( .A(pipeline_regfile_data[216]), .B(n13004), .S(n6650), .Z(
        n4820) );
  MUX2_X1 U7264 ( .A(pipeline_regfile_data[184]), .B(n9419), .S(n6651), .Z(
        n4819) );
  MUX2_X1 U7265 ( .A(pipeline_regfile_data[152]), .B(n13004), .S(n6652), .Z(
        n4818) );
  MUX2_X1 U7266 ( .A(pipeline_regfile_data[486]), .B(n9432), .S(n6644), .Z(
        n5387) );
  MUX2_X1 U7267 ( .A(pipeline_regfile_data[454]), .B(n13022), .S(n6645), .Z(
        n5386) );
  MUX2_X1 U7268 ( .A(pipeline_regfile_data[422]), .B(n9432), .S(n6646), .Z(
        n5385) );
  MUX2_X1 U7269 ( .A(pipeline_regfile_data[390]), .B(n13022), .S(n6647), .Z(
        n5384) );
  MUX2_X1 U7270 ( .A(pipeline_regfile_data[358]), .B(n9432), .S(n6648), .Z(
        n5383) );
  MUX2_X1 U7271 ( .A(pipeline_regfile_data[326]), .B(n13022), .S(n6653), .Z(
        n5382) );
  MUX2_X1 U7272 ( .A(pipeline_regfile_data[230]), .B(n9432), .S(n6649), .Z(
        n5379) );
  MUX2_X1 U7273 ( .A(pipeline_regfile_data[198]), .B(n13022), .S(n6650), .Z(
        n5378) );
  MUX2_X1 U7274 ( .A(pipeline_regfile_data[166]), .B(n9432), .S(n6651), .Z(
        n5377) );
  MUX2_X1 U7275 ( .A(pipeline_regfile_data[134]), .B(n13022), .S(n6652), .Z(
        n5376) );
  MUX2_X1 U7276 ( .A(pipeline_regfile_data[102]), .B(n9432), .S(n6654), .Z(
        n5375) );
  MUX2_X1 U7277 ( .A(pipeline_regfile_data[70]), .B(n13022), .S(n6655), .Z(
        n5374) );
  MUX2_X1 U7278 ( .A(pipeline_regfile_data[610]), .B(n9436), .S(n6671), .Z(
        n5515) );
  MUX2_X1 U7279 ( .A(pipeline_regfile_data[482]), .B(n9436), .S(n6644), .Z(
        n5511) );
  MUX2_X1 U7280 ( .A(pipeline_regfile_data[450]), .B(n13026), .S(n6645), .Z(
        n5510) );
  MUX2_X1 U7281 ( .A(pipeline_regfile_data[418]), .B(n9436), .S(n6646), .Z(
        n5509) );
  MUX2_X1 U7282 ( .A(pipeline_regfile_data[386]), .B(n13026), .S(n6647), .Z(
        n5508) );
  MUX2_X1 U7283 ( .A(pipeline_regfile_data[354]), .B(n9436), .S(n6648), .Z(
        n5507) );
  MUX2_X1 U7284 ( .A(pipeline_regfile_data[322]), .B(n13026), .S(n6653), .Z(
        n5506) );
  MUX2_X1 U7285 ( .A(pipeline_regfile_data[290]), .B(n9436), .S(n6656), .Z(
        n5505) );
  MUX2_X1 U7286 ( .A(pipeline_regfile_data[226]), .B(n9436), .S(n6649), .Z(
        n5503) );
  MUX2_X1 U7287 ( .A(pipeline_regfile_data[194]), .B(n13026), .S(n6650), .Z(
        n5502) );
  MUX2_X1 U7288 ( .A(pipeline_regfile_data[162]), .B(n9436), .S(n6651), .Z(
        n5501) );
  MUX2_X1 U7289 ( .A(pipeline_regfile_data[130]), .B(n13026), .S(n6652), .Z(
        n5500) );
  MUX2_X1 U7290 ( .A(pipeline_regfile_data[98]), .B(n9436), .S(n6654), .Z(
        n5499) );
  MUX2_X1 U7291 ( .A(pipeline_regfile_data[66]), .B(n13026), .S(n6655), .Z(
        n5498) );
  MUX2_X1 U7292 ( .A(pipeline_regfile_data[324]), .B(n13024), .S(n6653), .Z(
        n5444) );
  MUX2_X1 U7293 ( .A(pipeline_regfile_data[68]), .B(n13024), .S(n6655), .Z(
        n5436) );
  MUX2_X1 U7294 ( .A(pipeline_regfile_data[609]), .B(n9437), .S(n6671), .Z(
        n5546) );
  MUX2_X1 U7295 ( .A(pipeline_regfile_data[545]), .B(n9437), .S(n6672), .Z(
        n5544) );
  MUX2_X1 U7296 ( .A(pipeline_regfile_data[481]), .B(n9437), .S(n6644), .Z(
        n5542) );
  MUX2_X1 U7297 ( .A(pipeline_regfile_data[449]), .B(n13027), .S(n6645), .Z(
        n5541) );
  MUX2_X1 U7298 ( .A(pipeline_regfile_data[417]), .B(n9437), .S(n6646), .Z(
        n5540) );
  MUX2_X1 U7299 ( .A(pipeline_regfile_data[385]), .B(n13027), .S(n6647), .Z(
        n5539) );
  MUX2_X1 U7300 ( .A(pipeline_regfile_data[353]), .B(n9437), .S(n6648), .Z(
        n5538) );
  MUX2_X1 U7301 ( .A(pipeline_regfile_data[321]), .B(n13027), .S(n6653), .Z(
        n5537) );
  MUX2_X1 U7302 ( .A(pipeline_regfile_data[289]), .B(n9437), .S(n6656), .Z(
        n5536) );
  MUX2_X1 U7303 ( .A(pipeline_regfile_data[257]), .B(n13027), .S(n6657), .Z(
        n5535) );
  MUX2_X1 U7304 ( .A(pipeline_regfile_data[225]), .B(n9437), .S(n6649), .Z(
        n5534) );
  MUX2_X1 U7305 ( .A(pipeline_regfile_data[193]), .B(n13027), .S(n6650), .Z(
        n5533) );
  MUX2_X1 U7306 ( .A(pipeline_regfile_data[161]), .B(n9437), .S(n6651), .Z(
        n5532) );
  MUX2_X1 U7307 ( .A(pipeline_regfile_data[129]), .B(n13027), .S(n6652), .Z(
        n5531) );
  MUX2_X1 U7308 ( .A(pipeline_regfile_data[97]), .B(n9437), .S(n6654), .Z(
        n5530) );
  MUX2_X1 U7309 ( .A(pipeline_regfile_data[65]), .B(n13027), .S(n6655), .Z(
        n5529) );
  MUX2_X1 U7310 ( .A(pipeline_regfile_data[33]), .B(n9437), .S(n6658), .Z(
        n5528) );
  MUX2_X1 U7311 ( .A(pipeline_regfile_data[483]), .B(n9435), .S(n6644), .Z(
        n5480) );
  MUX2_X1 U7312 ( .A(pipeline_regfile_data[620]), .B(n9423), .S(n6671), .Z(
        n5205) );
  MUX2_X1 U7313 ( .A(pipeline_regfile_data[492]), .B(n9423), .S(n6644), .Z(
        n5201) );
  MUX2_X1 U7314 ( .A(pipeline_regfile_data[460]), .B(n13016), .S(n6645), .Z(
        n5200) );
  MUX2_X1 U7315 ( .A(pipeline_regfile_data[428]), .B(n9423), .S(n6646), .Z(
        n5199) );
  MUX2_X1 U7316 ( .A(pipeline_regfile_data[396]), .B(n13016), .S(n6647), .Z(
        n5198) );
  MUX2_X1 U7317 ( .A(pipeline_regfile_data[364]), .B(n9423), .S(n6648), .Z(
        n5197) );
  MUX2_X1 U7318 ( .A(pipeline_regfile_data[332]), .B(n13016), .S(n6653), .Z(
        n5196) );
  MUX2_X1 U7319 ( .A(pipeline_regfile_data[300]), .B(n9423), .S(n6656), .Z(
        n5195) );
  MUX2_X1 U7320 ( .A(pipeline_regfile_data[268]), .B(n13016), .S(n6657), .Z(
        n5194) );
  MUX2_X1 U7321 ( .A(pipeline_regfile_data[236]), .B(n9423), .S(n6649), .Z(
        n5193) );
  MUX2_X1 U7322 ( .A(pipeline_regfile_data[204]), .B(n13016), .S(n6650), .Z(
        n5192) );
  MUX2_X1 U7323 ( .A(pipeline_regfile_data[172]), .B(n9423), .S(n6651), .Z(
        n5191) );
  MUX2_X1 U7324 ( .A(pipeline_regfile_data[140]), .B(n13016), .S(n6652), .Z(
        n5190) );
  MUX2_X1 U7325 ( .A(pipeline_regfile_data[108]), .B(n9423), .S(n6654), .Z(
        n5189) );
  MUX2_X1 U7326 ( .A(pipeline_regfile_data[76]), .B(n13016), .S(n6655), .Z(
        n5188) );
  MUX2_X1 U7327 ( .A(pipeline_regfile_data[44]), .B(n9423), .S(n6658), .Z(
        n5187) );
  INV_X1 U7328 ( .A(pipeline_alu_src_b[26]), .ZN(n10016) );
  AND2_X1 U7329 ( .A1(pipeline_regfile_data[954]), .A2(n6728), .ZN(n7010) );
  AND2_X1 U7330 ( .A1(pipeline_regfile_data[698]), .A2(n6720), .ZN(n7011) );
  INV_X2 U7331 ( .A(n8244), .ZN(n8246) );
  INV_X2 U7332 ( .A(n8244), .ZN(n8247) );
  AND2_X1 U7333 ( .A1(n7012), .A2(n7013), .ZN(n7062) );
  NAND2_X1 U7334 ( .A1(n9925), .A2(n9924), .ZN(n7012) );
  NAND2_X1 U7335 ( .A1(n9928), .A2(n9927), .ZN(n7013) );
  INV_X2 U7336 ( .A(n9991), .ZN(n9817) );
  NAND2_X1 U7337 ( .A1(n7076), .A2(n10248), .ZN(n13099) );
  NAND2_X1 U7338 ( .A1(n9798), .A2(n9797), .ZN(n9915) );
  INV_X1 U7339 ( .A(n10056), .ZN(n9449) );
  NAND2_X1 U7341 ( .A1(n9705), .A2(n9797), .ZN(n9710) );
  INV_X4 U7342 ( .A(n9360), .ZN(imem_haddr[9]) );
  AND2_X4 U7343 ( .A1(n13097), .A2(n10258), .ZN(n7064) );
  OR2_X1 U7344 ( .A1(n11570), .A2(n12565), .ZN(n7066) );
  OR2_X1 U7345 ( .A1(n11414), .A2(n12565), .ZN(n7065) );
  OR2_X1 U7346 ( .A1(n11570), .A2(n9400), .ZN(n7067) );
  INV_X2 U7347 ( .A(n13105), .ZN(n11257) );
  INV_X2 U7348 ( .A(n13098), .ZN(n11105) );
  INV_X4 U7349 ( .A(n9630), .ZN(n7074) );
  INV_X4 U7350 ( .A(n6745), .ZN(n7073) );
  INV_X4 U7351 ( .A(n7072), .ZN(n9641) );
  AND2_X4 U7352 ( .A1(n7165), .A2(n10251), .ZN(n7077) );
  AND3_X1 U7353 ( .A1(n9648), .A2(n9650), .A3(pipeline_inst_DX[4]), .ZN(n7080)
         );
  NAND3_X1 U7354 ( .A1(n638), .A2(n637), .A3(n636), .ZN(n7014) );
  AND2_X1 U7355 ( .A1(n7054), .A2(n7163), .ZN(n7016) );
  AND3_X1 U7356 ( .A1(n12834), .A2(n6745), .A3(n9634), .ZN(n7083) );
  INV_X1 U7357 ( .A(n12394), .ZN(n12397) );
  AND3_X1 U7358 ( .A1(n6941), .A2(n12995), .A3(n12992), .ZN(n7087) );
  AND3_X1 U7359 ( .A1(n6941), .A2(n12996), .A3(n12992), .ZN(n7088) );
  NAND3_X1 U7360 ( .A1(n3785), .A2(n11741), .A3(n8223), .ZN(n11742) );
  NAND2_X1 U7361 ( .A1(n3785), .A2(n7167), .ZN(n10341) );
  NAND3_X1 U7362 ( .A1(n7054), .A2(n7078), .A3(n6843), .ZN(n10793) );
  AND3_X1 U7363 ( .A1(n693), .A2(pipeline_regfile_N18), .A3(n10336), .ZN(n7089) );
  AOI221_X1 U7364 ( .B1(pipeline_regfile_data[719]), .B2(n6734), .C1(
        pipeline_regfile_data[911]), .C2(n6733), .A(n7723), .ZN(n7698) );
  NOR4_X2 U7365 ( .A1(n7020), .A2(n7021), .A3(n7022), .A4(n7023), .ZN(n7122)
         );
  AOI221_X1 U7366 ( .B1(pipeline_regfile_data[735]), .B2(n6734), .C1(
        pipeline_regfile_data[927]), .C2(n6733), .A(n8237), .ZN(n8208) );
  AOI221_X1 U7367 ( .B1(pipeline_regfile_data[711]), .B2(n6734), .C1(
        pipeline_regfile_data[903]), .C2(n6733), .A(n7467), .ZN(n7442) );
  CLKBUF_X3 U7368 ( .A(n10339), .Z(n9402) );
  AOI221_X1 U7369 ( .B1(pipeline_regfile_data[704]), .B2(n6773), .C1(
        pipeline_regfile_data[896]), .C2(n6772), .A(n8303), .ZN(n8273) );
  AOI221_X1 U7370 ( .B1(pipeline_regfile_data[714]), .B2(n6734), .C1(
        pipeline_regfile_data[906]), .C2(n6733), .A(n7563), .ZN(n7538) );
  AOI221_X1 U7371 ( .B1(pipeline_regfile_data[718]), .B2(n6734), .C1(
        pipeline_regfile_data[910]), .C2(n6733), .A(n7691), .ZN(n7666) );
  AOI221_X1 U7372 ( .B1(pipeline_regfile_data[735]), .B2(n6773), .C1(
        pipeline_regfile_data[927]), .C2(n6772), .A(n9295), .ZN(n9264) );
  AOI221_X1 U7373 ( .B1(pipeline_regfile_data[710]), .B2(n6734), .C1(
        pipeline_regfile_data[902]), .C2(n6733), .A(n7435), .ZN(n7410) );
  AOI221_X1 U7374 ( .B1(pipeline_regfile_data[719]), .B2(n6773), .C1(
        pipeline_regfile_data[911]), .C2(n6772), .A(n8779), .ZN(n8754) );
  AOI221_X1 U7375 ( .B1(pipeline_regfile_data[535]), .B2(n6709), .C1(
        pipeline_regfile_data[983]), .C2(n6763), .A(n9036), .ZN(n9007) );
  AOI221_X1 U7376 ( .B1(pipeline_regfile_data[725]), .B2(n6773), .C1(
        pipeline_regfile_data[917]), .C2(n6772), .A(n8971), .ZN(n8946) );
  AOI221_X1 U7377 ( .B1(pipeline_regfile_data[729]), .B2(n6773), .C1(
        pipeline_regfile_data[921]), .C2(n6772), .A(n9097), .ZN(n9072) );
  AOI221_X1 U7378 ( .B1(pipeline_regfile_data[722]), .B2(n6773), .C1(
        pipeline_regfile_data[914]), .C2(n6772), .A(n8875), .ZN(n8850) );
  AOI221_X1 U7379 ( .B1(pipeline_regfile_data[728]), .B2(n6773), .C1(
        pipeline_regfile_data[920]), .C2(n6772), .A(n9065), .ZN(n9040) );
  AOI221_X1 U7380 ( .B1(pipeline_regfile_data[721]), .B2(n6773), .C1(
        pipeline_regfile_data[913]), .C2(n6772), .A(n8843), .ZN(n8818) );
  AOI221_X1 U7381 ( .B1(pipeline_regfile_data[724]), .B2(n6773), .C1(
        pipeline_regfile_data[916]), .C2(n6772), .A(n8939), .ZN(n8914) );
  AOI221_X1 U7382 ( .B1(pipeline_regfile_data[726]), .B2(n6773), .C1(
        pipeline_regfile_data[918]), .C2(n6772), .A(n9001), .ZN(n8978) );
  AOI221_X1 U7383 ( .B1(pipeline_regfile_data[723]), .B2(n6773), .C1(
        pipeline_regfile_data[915]), .C2(n6772), .A(n8907), .ZN(n8882) );
  AOI221_X1 U7384 ( .B1(pipeline_regfile_data[734]), .B2(n6773), .C1(
        pipeline_regfile_data[926]), .C2(n6772), .A(n9257), .ZN(n9232) );
  AOI221_X1 U7385 ( .B1(pipeline_regfile_data[733]), .B2(n6773), .C1(
        pipeline_regfile_data[925]), .C2(n6772), .A(n9225), .ZN(n9200) );
  AOI221_X1 U7386 ( .B1(pipeline_regfile_data[730]), .B2(n6773), .C1(
        pipeline_regfile_data[922]), .C2(n6772), .A(n9129), .ZN(n9104) );
  AOI221_X1 U7387 ( .B1(pipeline_regfile_data[732]), .B2(n6773), .C1(
        pipeline_regfile_data[924]), .C2(n6772), .A(n9193), .ZN(n9168) );
  AOI221_X1 U7388 ( .B1(pipeline_regfile_data[717]), .B2(n6734), .C1(
        pipeline_regfile_data[909]), .C2(n6733), .A(n7659), .ZN(n7634) );
  AOI221_X1 U7389 ( .B1(pipeline_regfile_data[709]), .B2(n6734), .C1(
        pipeline_regfile_data[901]), .C2(n6733), .A(n7403), .ZN(n7378) );
  AOI221_X1 U7390 ( .B1(pipeline_regfile_data[713]), .B2(n6734), .C1(
        pipeline_regfile_data[905]), .C2(n6733), .A(n7531), .ZN(n7506) );
  AOI221_X1 U7391 ( .B1(pipeline_regfile_data[714]), .B2(n6773), .C1(
        pipeline_regfile_data[906]), .C2(n6772), .A(n8619), .ZN(n8594) );
  AOI221_X1 U7392 ( .B1(pipeline_regfile_data[729]), .B2(n6734), .C1(
        pipeline_regfile_data[921]), .C2(n6733), .A(n8042), .ZN(n8017) );
  AOI221_X1 U7393 ( .B1(pipeline_regfile_data[727]), .B2(n6734), .C1(
        pipeline_regfile_data[919]), .C2(n6733), .A(n7978), .ZN(n7953) );
  AOI221_X1 U7394 ( .B1(pipeline_regfile_data[731]), .B2(n6734), .C1(
        pipeline_regfile_data[923]), .C2(n6733), .A(n8105), .ZN(n8080) );
  NOR4_X2 U7395 ( .A1(n7027), .A2(n7028), .A3(n7029), .A4(n7030), .ZN(n7127)
         );
  NOR4_X2 U7396 ( .A1(n7031), .A2(n7032), .A3(n7033), .A4(n7034), .ZN(n7128)
         );
  AOI221_X1 U7397 ( .B1(pipeline_regfile_data[725]), .B2(n6734), .C1(
        pipeline_regfile_data[917]), .C2(n6733), .A(n7914), .ZN(n7889) );
  NOR4_X2 U7398 ( .A1(n7035), .A2(n7036), .A3(n7037), .A4(n6785), .ZN(n7130)
         );
  AOI221_X1 U7399 ( .B1(pipeline_regfile_data[720]), .B2(n6734), .C1(
        pipeline_regfile_data[912]), .C2(n6733), .A(n7755), .ZN(n7730) );
  AOI221_X1 U7400 ( .B1(pipeline_regfile_data[722]), .B2(n6734), .C1(
        pipeline_regfile_data[914]), .C2(n6733), .A(n7818), .ZN(n7793) );
  AOI221_X1 U7401 ( .B1(pipeline_regfile_data[723]), .B2(n6734), .C1(
        pipeline_regfile_data[915]), .C2(n6733), .A(n7850), .ZN(n7825) );
  AOI221_X1 U7402 ( .B1(pipeline_regfile_data[726]), .B2(n6734), .C1(
        pipeline_regfile_data[918]), .C2(n6733), .A(n7946), .ZN(n7921) );
  AOI221_X1 U7403 ( .B1(pipeline_regfile_data[732]), .B2(n6734), .C1(
        pipeline_regfile_data[924]), .C2(n6733), .A(n8137), .ZN(n8112) );
  AOI221_X1 U7404 ( .B1(pipeline_regfile_data[733]), .B2(n6734), .C1(
        pipeline_regfile_data[925]), .C2(n6733), .A(n8169), .ZN(n8144) );
  AOI221_X1 U7405 ( .B1(pipeline_regfile_data[712]), .B2(n6734), .C1(
        pipeline_regfile_data[904]), .C2(n6733), .A(n7499), .ZN(n7474) );
  AOI221_X1 U7406 ( .B1(pipeline_regfile_data[712]), .B2(n6773), .C1(
        pipeline_regfile_data[904]), .C2(n6772), .A(n8555), .ZN(n8530) );
  AOI221_X1 U7407 ( .B1(pipeline_regfile_data[716]), .B2(n6773), .C1(
        pipeline_regfile_data[908]), .C2(n6772), .A(n8683), .ZN(n8658) );
  NOR4_X2 U7408 ( .A1(n7046), .A2(n7047), .A3(n7048), .A4(n7049), .ZN(n7144)
         );
  AOI221_X1 U7409 ( .B1(pipeline_regfile_data[715]), .B2(n6773), .C1(
        pipeline_regfile_data[907]), .C2(n6772), .A(n8651), .ZN(n8626) );
  AOI221_X1 U7410 ( .B1(pipeline_regfile_data[709]), .B2(n6773), .C1(
        pipeline_regfile_data[901]), .C2(n6772), .A(n8459), .ZN(n8434) );
  NOR2_X1 U7411 ( .A1(n12462), .A2(n9485), .ZN(n12463) );
  INV_X4 U7412 ( .A(n9079), .ZN(n7156) );
  INV_X4 U7413 ( .A(n9078), .ZN(n7155) );
  INV_X4 U7414 ( .A(n8633), .ZN(n7158) );
  INV_X4 U7415 ( .A(n8632), .ZN(n7157) );
  INV_X4 U7416 ( .A(n8697), .ZN(n7160) );
  INV_X4 U7417 ( .A(n8696), .ZN(n7159) );
  INV_X4 U7418 ( .A(n9142), .ZN(n7149) );
  OAI22_X1 U7419 ( .A1(n6639), .A2(n10126), .B1(n693), .B2(n12823), .ZN(n6283)
         );
  AND2_X4 U7420 ( .A1(n7075), .A2(n702), .ZN(n7165) );
  AOI221_X1 U7421 ( .B1(pipeline_regfile_data[713]), .B2(n6773), .C1(
        pipeline_regfile_data[905]), .C2(n6772), .A(n8587), .ZN(n8562) );
  AND3_X1 U7422 ( .A1(pipeline_inst_DX[30]), .A2(n10242), .A3(n7055), .ZN(
        n7163) );
  AND2_X4 U7423 ( .A1(pipeline_regfile_N19), .A2(n7078), .ZN(n7169) );
  AND3_X1 U7424 ( .A1(n9632), .A2(n8223), .A3(n9617), .ZN(n7182) );
  AND2_X4 U7425 ( .A1(n7165), .A2(n8214), .ZN(n7176) );
  AND2_X2 U7426 ( .A1(n10336), .A2(n8214), .ZN(n7172) );
  INV_X4 U7427 ( .A(n9015), .ZN(n7152) );
  INV_X4 U7428 ( .A(n9014), .ZN(n7151) );
  INV_X4 U7429 ( .A(n8953), .ZN(n7154) );
  INV_X4 U7430 ( .A(n8952), .ZN(n7153) );
  INV_X4 U7431 ( .A(n8793), .ZN(n7162) );
  INV_X4 U7432 ( .A(n8792), .ZN(n7161) );
  AND3_X1 U7433 ( .A1(dmem_hsize[1]), .A2(n13096), .A3(n7064), .ZN(n7168) );
  AND2_X1 U7434 ( .A1(n7174), .A2(n693), .ZN(n7051) );
  XNOR2_X1 U7435 ( .A(pipeline_regfile_N15), .B(n12995), .ZN(n9646) );
  AND2_X4 U7436 ( .A1(n9631), .A2(pipeline_inst_DX[5]), .ZN(n7173) );
  NAND2_X1 U7437 ( .A1(n9721), .A2(n9651), .ZN(n7052) );
  NAND3_X1 U7438 ( .A1(pipeline_regfile_N12), .A2(n638), .A3(n637), .ZN(n7053)
         );
  AND3_X2 U7439 ( .A1(n10236), .A2(n10235), .A3(n10336), .ZN(n7054) );
  AND2_X1 U7440 ( .A1(pipeline_inst_DX[29]), .A2(pipeline_inst_DX[28]), .ZN(
        n7055) );
  AND2_X1 U7441 ( .A1(n6795), .A2(n601), .ZN(n7184) );
  AOI221_X1 U7442 ( .B1(pipeline_csr_mtvec[5]), .B2(n11229), .C1(
        pipeline_csr_mtime_full[37]), .C2(n9528), .A(n10782), .ZN(n10789) );
  OAI22_X1 U7443 ( .A1(n13111), .A2(n6901), .B1(n11269), .B2(n10947), .ZN(
        n10948) );
  OAI22_X1 U7444 ( .A1(n13111), .A2(n6902), .B1(n11269), .B2(n11054), .ZN(
        n11055) );
  OAI22_X1 U7445 ( .A1(n13111), .A2(n6903), .B1(n11269), .B2(n11081), .ZN(
        n11082) );
  OAI22_X1 U7446 ( .A1(n13111), .A2(n6904), .B1(n11269), .B2(n11139), .ZN(
        n11140) );
  OAI22_X1 U7447 ( .A1(n13111), .A2(n6905), .B1(n11269), .B2(n11027), .ZN(
        n11028) );
  OAI22_X1 U7448 ( .A1(n13111), .A2(n6906), .B1(n11269), .B2(n10866), .ZN(
        n10867) );
  OAI22_X1 U7449 ( .A1(n13111), .A2(n6907), .B1(n11269), .B2(n10920), .ZN(
        n10921) );
  OAI22_X1 U7450 ( .A1(n13111), .A2(n6908), .B1(n11269), .B2(n10974), .ZN(
        n10975) );
  OAI22_X1 U7451 ( .A1(n13111), .A2(n6909), .B1(n11269), .B2(n10839), .ZN(
        n10840) );
  OAI22_X1 U7452 ( .A1(n13111), .A2(n6910), .B1(n11269), .B2(n10754), .ZN(
        n10755) );
  OAI22_X1 U7453 ( .A1(n13111), .A2(n6911), .B1(n11269), .B2(n10243), .ZN(
        n10244) );
  NOR2_X1 U7454 ( .A1(pipeline_regfile_N18), .A2(n10333), .ZN(n10334) );
  AND2_X4 U7455 ( .A1(n6941), .A2(n12993), .ZN(n7191) );
  AND3_X1 U7456 ( .A1(pipeline_regfile_N17), .A2(n6628), .A3(n7181), .ZN(n7192) );
  MUX2_X1 U7457 ( .A(pipeline_regfile_data[507]), .B(n9416), .S(n6644), .Z(
        n4736) );
  MUX2_X1 U7458 ( .A(pipeline_regfile_data[443]), .B(n9416), .S(n6646), .Z(
        n4734) );
  MUX2_X1 U7459 ( .A(pipeline_regfile_data[379]), .B(n9416), .S(n6648), .Z(
        n4732) );
  MUX2_X1 U7460 ( .A(pipeline_regfile_data[475]), .B(n13001), .S(n6645), .Z(
        n4735) );
  MUX2_X1 U7461 ( .A(pipeline_regfile_data[411]), .B(n13001), .S(n6647), .Z(
        n4733) );
  MUX2_X1 U7462 ( .A(pipeline_regfile_data[491]), .B(n9425), .S(n6644), .Z(
        n5232) );
  MUX2_X1 U7463 ( .A(pipeline_regfile_data[459]), .B(n13017), .S(n6645), .Z(
        n5231) );
  MUX2_X1 U7464 ( .A(pipeline_regfile_data[427]), .B(n9424), .S(n6646), .Z(
        n5230) );
  MUX2_X1 U7465 ( .A(pipeline_regfile_data[395]), .B(n9425), .S(n6647), .Z(
        n5229) );
  MUX2_X1 U7466 ( .A(pipeline_regfile_data[356]), .B(n9434), .S(n6648), .Z(
        n5445) );
  MUX2_X1 U7467 ( .A(pipeline_regfile_data[100]), .B(n9434), .S(n6654), .Z(
        n5437) );
  MUX2_X1 U7468 ( .A(pipeline_regfile_data[493]), .B(n9422), .S(n6644), .Z(
        n5170) );
  MUX2_X1 U7469 ( .A(pipeline_regfile_data[461]), .B(n13015), .S(n6645), .Z(
        n5169) );
  MUX2_X1 U7470 ( .A(pipeline_regfile_data[429]), .B(n9422), .S(n6646), .Z(
        n5168) );
  MUX2_X1 U7471 ( .A(pipeline_regfile_data[397]), .B(n13015), .S(n6647), .Z(
        n5167) );
  AOI221_X1 U7472 ( .B1(pipeline_csr_time_full[6]), .B2(n6735), .C1(
        pipeline_csr_cycle_full[6]), .C2(n13116), .A(n10734), .ZN(n10735) );
  AOI221_X1 U7473 ( .B1(pipeline_csr_mtime_full[60]), .B2(n9528), .C1(
        pipeline_csr_from_host[28]), .C2(n9461), .A(n10432), .ZN(n10436) );
  AOI221_X1 U7474 ( .B1(pipeline_csr_time_full[20]), .B2(n6735), .C1(
        pipeline_csr_cycle_full[20]), .C2(n13116), .A(n10894), .ZN(n10903) );
  AOI221_X1 U7475 ( .B1(pipeline_csr_time_full[15]), .B2(n6735), .C1(
        pipeline_csr_cycle_full[15]), .C2(n13116), .A(n11110), .ZN(n11120) );
  AOI221_X1 U7476 ( .B1(pipeline_csr_time_full[8]), .B2(n6735), .C1(
        pipeline_csr_cycle_full[8]), .C2(n13116), .A(n10623), .ZN(n10630) );
  AND2_X1 U7477 ( .A1(pipeline_ctrl_prev_ex_code_WB[1]), .A2(
        pipeline_ctrl_had_ex_WB), .ZN(n7216) );
  NAND3_X1 U7478 ( .A1(n7163), .A2(n693), .A3(n6847), .ZN(n10825) );
  AOI221_X1 U7479 ( .B1(pipeline_md_N32), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[3]), .A(n10480), .ZN(n10481) );
  NAND2_X1 U7480 ( .A1(n603), .A2(pipeline_rs1_data_bypassed[3]), .ZN(n10502)
         );
  NAND2_X2 U7481 ( .A1(pipeline_alu_N90), .A2(n6813), .ZN(n7058) );
  INV_X4 U7482 ( .A(n12594), .ZN(n7060) );
  INV_X4 U7483 ( .A(n6643), .ZN(n9521) );
  INV_X4 U7484 ( .A(n12827), .ZN(n9524) );
  INV_X4 U7485 ( .A(n12827), .ZN(n9523) );
  INV_X4 U7486 ( .A(n12827), .ZN(n9525) );
  INV_X4 U7487 ( .A(n9458), .ZN(n9454) );
  INV_X4 U7488 ( .A(n6777), .ZN(n9497) );
  INV_X4 U7489 ( .A(n6777), .ZN(n9496) );
  INV_X4 U7490 ( .A(n9458), .ZN(n9455) );
  INV_X4 U7491 ( .A(n6573), .ZN(n9458) );
  INV_X4 U7492 ( .A(n9457), .ZN(n9456) );
  INV_X4 U7493 ( .A(n9459), .ZN(n9453) );
  INV_X4 U7494 ( .A(n9452), .ZN(n9450) );
  INV_X4 U7495 ( .A(n9452), .ZN(n9451) );
  INV_X4 U7496 ( .A(n9513), .ZN(n9512) );
  INV_X4 U7497 ( .A(n9508), .ZN(n9507) );
  INV_X4 U7498 ( .A(n9506), .ZN(n9505) );
  INV_X4 U7499 ( .A(n6643), .ZN(n9520) );
  INV_X4 U7500 ( .A(n9473), .ZN(n9472) );
  AOI22_X1 U7501 ( .A1(n9977), .A2(n9818), .B1(n9989), .B2(n9817), .ZN(n9996)
         );
  AOI22_X1 U7502 ( .A1(n10007), .A2(n9810), .B1(n10018), .B2(n9809), .ZN(
        n10025) );
  AOI22_X2 U7503 ( .A1(n10035), .A2(n9804), .B1(n10047), .B2(n9803), .ZN(
        n10054) );
  AOI22_X2 U7504 ( .A1(n10039), .A2(n10038), .B1(n10037), .B2(n10036), .ZN(
        n10040) );
  OAI211_X2 U7505 ( .C1(n7062), .C2(n9938), .A(n9937), .B(n9936), .ZN(n9952)
         );
  NAND2_X2 U7506 ( .A1(n9873), .A2(n9888), .ZN(n9882) );
  INV_X4 U7507 ( .A(n12565), .ZN(n9489) );
  INV_X4 U7508 ( .A(n6780), .ZN(n9487) );
  INV_X4 U7509 ( .A(n9444), .ZN(n9443) );
  INV_X4 U7510 ( .A(n7014), .ZN(n9326) );
  INV_X4 U7511 ( .A(n7014), .ZN(n9327) );
  INV_X4 U7512 ( .A(n11261), .ZN(n9527) );
  NAND2_X2 U7513 ( .A1(n12411), .A2(n12412), .ZN(n12556) );
  INV_X4 U7514 ( .A(n9307), .ZN(n9309) );
  INV_X4 U7515 ( .A(n9307), .ZN(n9310) );
  INV_X4 U7516 ( .A(n11574), .ZN(n9471) );
  INV_X4 U7517 ( .A(n12645), .ZN(n9511) );
  INV_X4 U7518 ( .A(n10276), .ZN(n9500) );
  INV_X4 U7519 ( .A(n10276), .ZN(n9499) );
  INV_X4 U7520 ( .A(n9510), .ZN(n9509) );
  INV_X4 U7521 ( .A(n12687), .ZN(n12749) );
  AOI21_X2 U7522 ( .B1(n12305), .B2(n9511), .A(n11686), .ZN(n11725) );
  AOI21_X2 U7523 ( .B1(n12642), .B2(n9511), .A(n11769), .ZN(n11802) );
  AOI21_X2 U7524 ( .B1(n12576), .B2(n9511), .A(n11841), .ZN(n11878) );
  INV_X4 U7525 ( .A(n12783), .ZN(n9513) );
  INV_X4 U7526 ( .A(n12765), .ZN(n9506) );
  INV_X4 U7527 ( .A(n12774), .ZN(n9508) );
  NAND2_X2 U7528 ( .A1(n12172), .A2(n9510), .ZN(n12182) );
  INV_X4 U7529 ( .A(n12785), .ZN(n12172) );
  INV_X4 U7530 ( .A(n12763), .ZN(n9503) );
  INV_X4 U7531 ( .A(n13099), .ZN(n11233) );
  INV_X4 U7532 ( .A(n12346), .ZN(n9473) );
  INV_X4 U7533 ( .A(n9477), .ZN(n9476) );
  INV_X4 U7534 ( .A(n12347), .ZN(n9474) );
  AOI21_X2 U7535 ( .B1(n9490), .B2(n9468), .A(n10516), .ZN(n9404) );
  AOI21_X2 U7536 ( .B1(n9490), .B2(n9468), .A(n10516), .ZN(n12257) );
  INV_X4 U7537 ( .A(n11283), .ZN(n9468) );
  INV_X4 U7538 ( .A(n12827), .ZN(n9522) );
  INV_X4 U7539 ( .A(n6640), .ZN(n9460) );
  INV_X4 U7540 ( .A(n9514), .ZN(n9515) );
  INV_X4 U7541 ( .A(n6706), .ZN(n9529) );
  INV_X4 U7542 ( .A(n11572), .ZN(n12276) );
  INV_X4 U7543 ( .A(n12273), .ZN(n11869) );
  INV_X4 U7544 ( .A(n9785), .ZN(n9444) );
  INV_X4 U7545 ( .A(n8245), .ZN(n8244) );
  INV_X4 U7546 ( .A(n9311), .ZN(n9307) );
  INV_X8 U7547 ( .A(n9364), .ZN(imem_haddr[25]) );
  AND2_X1 U7548 ( .A1(n10248), .A2(n10251), .ZN(n7063) );
  INV_X4 U7549 ( .A(n9495), .ZN(n9494) );
  INV_X4 U7550 ( .A(n6737), .ZN(n9493) );
  INV_X4 U7551 ( .A(n6735), .ZN(n9526) );
  INV_X4 U7552 ( .A(n9312), .ZN(n9315) );
  INV_X4 U7553 ( .A(n9312), .ZN(n9316) );
  INV_X4 U7554 ( .A(n9449), .ZN(n9448) );
  INV_X4 U7555 ( .A(n9322), .ZN(n9325) );
  INV_X4 U7556 ( .A(n7050), .ZN(n8270) );
  INV_X4 U7557 ( .A(n6580), .ZN(n8266) );
  INV_X4 U7558 ( .A(n9317), .ZN(n9319) );
  INV_X4 U7559 ( .A(n6696), .ZN(n8256) );
  INV_X4 U7560 ( .A(n6580), .ZN(n8268) );
  INV_X4 U7561 ( .A(n7050), .ZN(n8269) );
  INV_X4 U7562 ( .A(n6696), .ZN(n8255) );
  AND2_X1 U7563 ( .A1(n11690), .A2(n7065), .ZN(n11332) );
  AND2_X1 U7564 ( .A1(n11618), .A2(n7066), .ZN(n11156) );
  INV_X4 U7565 ( .A(n12776), .ZN(n9510) );
  INV_X4 U7566 ( .A(n6665), .ZN(n9463) );
  INV_X4 U7567 ( .A(n6666), .ZN(n9467) );
  NAND2_X2 U7568 ( .A1(n12662), .A2(n12800), .ZN(n12785) );
  INV_X4 U7569 ( .A(n12355), .ZN(n12793) );
  AND2_X1 U7570 ( .A1(n11569), .A2(n7067), .ZN(n11571) );
  INV_X4 U7571 ( .A(n9502), .ZN(n9501) );
  NAND2_X2 U7573 ( .A1(n12567), .A2(n12800), .ZN(n12639) );
  NAND2_X2 U7574 ( .A1(n11159), .A2(n12800), .ZN(n12772) );
  AND2_X1 U7575 ( .A1(n10082), .A2(n9800), .ZN(n7068) );
  INV_X4 U7576 ( .A(n12357), .ZN(n9479) );
  INV_X4 U7577 ( .A(n13113), .ZN(n11268) );
  AOI21_X2 U7578 ( .B1(n9491), .B2(n9468), .A(n11198), .ZN(n11284) );
  INV_X4 U7579 ( .A(n12350), .ZN(n9477) );
  INV_X4 U7580 ( .A(n6697), .ZN(n9462) );
  AND2_X1 U7581 ( .A1(n10082), .A2(n10081), .ZN(n7069) );
  INV_X4 U7582 ( .A(n9491), .ZN(n9492) );
  AOI21_X2 U7583 ( .B1(n9470), .B2(n9468), .A(n10516), .ZN(n9405) );
  AOI21_X2 U7584 ( .B1(n9470), .B2(n9468), .A(n10516), .ZN(n9406) );
  INV_X4 U7585 ( .A(n12617), .ZN(n12809) );
  INV_X4 U7586 ( .A(n13104), .ZN(n11229) );
  INV_X4 U7587 ( .A(n13103), .ZN(n11136) );
  INV_X4 U7588 ( .A(n13114), .ZN(n11138) );
  INV_X4 U7589 ( .A(n12612), .ZN(n9490) );
  INV_X4 U7590 ( .A(n12892), .ZN(n12983) );
  INV_X4 U7591 ( .A(n12349), .ZN(n9475) );
  INV_X4 U7592 ( .A(n6670), .ZN(n9498) );
  INV_X4 U7593 ( .A(n9470), .ZN(n9469) );
  INV_X4 U7594 ( .A(n6849), .ZN(n9516) );
  INV_X4 U7595 ( .A(n9531), .ZN(n9530) );
  INV_X4 U7596 ( .A(n12899), .ZN(n12896) );
  NAND2_X2 U7597 ( .A1(n7076), .A2(n7051), .ZN(n13098) );
  INV_X4 U7598 ( .A(n8278), .ZN(n9304) );
  NAND2_X2 U7599 ( .A1(n7076), .A2(n7165), .ZN(n13105) );
  NAND2_X2 U7600 ( .A1(n7163), .A2(n7077), .ZN(n11264) );
  NAND2_X2 U7601 ( .A1(n7166), .A2(n7165), .ZN(n13114) );
  INV_X4 U7602 ( .A(n12839), .ZN(n9781) );
  NAND2_X2 U7603 ( .A1(n9820), .A2(pipeline_imm_31_), .ZN(n10043) );
  AND2_X1 U7604 ( .A1(n10333), .A2(n9658), .ZN(n7075) );
  INV_X4 U7605 ( .A(n11235), .ZN(n9461) );
  INV_X4 U7606 ( .A(n12632), .ZN(n9495) );
  AND2_X1 U7607 ( .A1(n7079), .A2(n9402), .ZN(n7076) );
  INV_X4 U7608 ( .A(pipeline_rs1_data_bypassed[3]), .ZN(n12526) );
  INV_X4 U7609 ( .A(n9318), .ZN(n9317) );
  INV_X4 U7610 ( .A(n7226), .ZN(n8250) );
  INV_X4 U7611 ( .A(n8285), .ZN(n9322) );
  INV_X4 U7612 ( .A(n11269), .ZN(n9466) );
  AND2_X1 U7613 ( .A1(n6796), .A2(n7172), .ZN(n7079) );
  INV_X4 U7614 ( .A(n9535), .ZN(n9534) );
  AND2_X1 U7615 ( .A1(n6641), .A2(n10251), .ZN(n7081) );
  AND4_X2 U7616 ( .A1(n11873), .A2(n11872), .A3(n11871), .A4(n11870), .ZN(
        n7082) );
  INV_X4 U7617 ( .A(n10416), .ZN(n1909) );
  INV_X4 U7618 ( .A(n11892), .ZN(n11943) );
  INV_X4 U7619 ( .A(n10422), .ZN(n12601) );
  AND3_X2 U7620 ( .A1(n9489), .A2(n9399), .A3(pipeline_alu_src_a[0]), .ZN(
        n7084) );
  NAND2_X2 U7621 ( .A1(n10085), .A2(n10083), .ZN(n12355) );
  AND3_X2 U7622 ( .A1(n9643), .A2(n7086), .A3(n6664), .ZN(n7085) );
  INV_X4 U7623 ( .A(n11739), .ZN(n11752) );
  INV_X4 U7624 ( .A(n12753), .ZN(n9502) );
  AND3_X2 U7625 ( .A1(n10242), .A2(n9634), .A3(n9633), .ZN(n7086) );
  NAND2_X2 U7626 ( .A1(n12062), .A2(n7005), .ZN(n12659) );
  INV_X4 U7627 ( .A(n12823), .ZN(n9517) );
  OAI221_X2 U7628 ( .B1(n12852), .B2(n9407), .C1(n9409), .C2(n12851), .A(
        n12865), .ZN(n9412) );
  OAI221_X2 U7629 ( .B1(n12854), .B2(n9407), .C1(n12892), .C2(n12853), .A(
        n12865), .ZN(n9413) );
  OAI221_X2 U7630 ( .B1(n12856), .B2(n9407), .C1(n9408), .C2(n12855), .A(
        n12865), .ZN(n9414) );
  OAI221_X2 U7631 ( .B1(n12858), .B2(n9407), .C1(n9409), .C2(n12857), .A(
        n12865), .ZN(n9415) );
  OAI221_X1 U7632 ( .B1(n12860), .B2(n9407), .C1(n12892), .C2(n12859), .A(
        n12865), .ZN(n9416) );
  OAI221_X2 U7633 ( .B1(n12862), .B2(n9407), .C1(n9408), .C2(n12861), .A(
        n12865), .ZN(n9417) );
  OAI221_X2 U7634 ( .B1(n12864), .B2(n9407), .C1(n9409), .C2(n12863), .A(
        n12865), .ZN(n9418) );
  OAI221_X2 U7635 ( .B1(n12867), .B2(n9407), .C1(n12892), .C2(n12866), .A(
        n12865), .ZN(n9419) );
  OAI221_X2 U7636 ( .B1(n12852), .B2(n9407), .C1(n9408), .C2(n12851), .A(
        n12865), .ZN(n12997) );
  OAI221_X2 U7637 ( .B1(n12854), .B2(n9407), .C1(n9409), .C2(n12853), .A(
        n12865), .ZN(n12998) );
  OAI221_X2 U7638 ( .B1(n12856), .B2(n9407), .C1(n12892), .C2(n12855), .A(
        n12865), .ZN(n12999) );
  OAI221_X2 U7639 ( .B1(n12858), .B2(n9407), .C1(n9408), .C2(n12857), .A(
        n12865), .ZN(n13000) );
  OAI221_X1 U7640 ( .B1(n12860), .B2(n9407), .C1(n9409), .C2(n12859), .A(
        n12865), .ZN(n13001) );
  OAI221_X2 U7641 ( .B1(n12862), .B2(n9407), .C1(n12892), .C2(n12861), .A(
        n12865), .ZN(n13002) );
  OAI221_X2 U7642 ( .B1(n12864), .B2(n9407), .C1(n9408), .C2(n12863), .A(
        n12865), .ZN(n13003) );
  OAI221_X2 U7643 ( .B1(n12867), .B2(n9407), .C1(n9409), .C2(n12866), .A(
        n12865), .ZN(n13004) );
  NAND2_X2 U7644 ( .A1(n12936), .A2(n12937), .ZN(n12892) );
  NAND4_X2 U7645 ( .A1(n12849), .A2(n12848), .A3(n12847), .A4(n12846), .ZN(
        n12940) );
  INV_X4 U7647 ( .A(n12352), .ZN(n9478) );
  INV_X4 U7648 ( .A(n12258), .ZN(n9470) );
  OAI221_X2 U7649 ( .B1(n12904), .B2(n9407), .C1(n12903), .C2(n12902), .A(
        n9410), .ZN(n9420) );
  OAI221_X2 U7650 ( .B1(n12910), .B2(n12909), .C1(n12908), .C2(n9407), .A(
        n12940), .ZN(n9421) );
  OAI221_X2 U7651 ( .B1(n12915), .B2(n12914), .C1(n12913), .C2(n9407), .A(
        n9411), .ZN(n9422) );
  OAI221_X2 U7652 ( .B1(n12920), .B2(n12919), .C1(n12918), .C2(n9407), .A(
        n9410), .ZN(n9423) );
  OAI221_X2 U7653 ( .B1(n12904), .B2(n9407), .C1(n12903), .C2(n12902), .A(
        n9411), .ZN(n13013) );
  OAI221_X2 U7654 ( .B1(n12910), .B2(n12909), .C1(n12908), .C2(n9407), .A(
        n9410), .ZN(n13014) );
  OAI221_X2 U7655 ( .B1(n12915), .B2(n12914), .C1(n12913), .C2(n9407), .A(
        n12940), .ZN(n13015) );
  OAI221_X2 U7656 ( .B1(n12920), .B2(n12919), .C1(n12918), .C2(n9407), .A(
        n9411), .ZN(n13016) );
  NAND2_X2 U7657 ( .A1(n12936), .A2(n12937), .ZN(n9408) );
  NAND2_X2 U7658 ( .A1(n12936), .A2(n12937), .ZN(n9409) );
  NAND4_X2 U7659 ( .A1(n12849), .A2(n12848), .A3(n12847), .A4(n12846), .ZN(
        n9410) );
  NAND4_X2 U7660 ( .A1(n12849), .A2(n12848), .A3(n12847), .A4(n12846), .ZN(
        n9411) );
  INV_X4 U7661 ( .A(n12806), .ZN(n12668) );
  INV_X4 U7662 ( .A(n3704), .ZN(n13131) );
  INV_X8 U7663 ( .A(n12945), .ZN(n9407) );
  INV_X4 U7664 ( .A(n3689), .ZN(n9531) );
  INV_X4 U7665 ( .A(n4231), .ZN(n13144) );
  AND4_X2 U7666 ( .A1(n8785), .A2(n8786), .A3(n8787), .A4(n8788), .ZN(n7091)
         );
  AND4_X2 U7667 ( .A1(n8272), .A2(n8273), .A3(n8274), .A4(n8275), .ZN(n7093)
         );
  AND4_X2 U7668 ( .A1(n7537), .A2(n7538), .A3(n7539), .A4(n7540), .ZN(n7094)
         );
  AND4_X2 U7669 ( .A1(n7409), .A2(n7410), .A3(n7411), .A4(n7412), .ZN(n7098)
         );
  AND4_X2 U7670 ( .A1(n7697), .A2(n7698), .A3(n7699), .A4(n7700), .ZN(n7100)
         );
  AND4_X2 U7671 ( .A1(n8497), .A2(n8498), .A3(n8499), .A4(n8500), .ZN(n7104)
         );
  AND4_X2 U7672 ( .A1(n9039), .A2(n9040), .A3(n9041), .A4(n9042), .ZN(n7107)
         );
  AND4_X2 U7673 ( .A1(n8817), .A2(n8818), .A3(n8819), .A4(n8820), .ZN(n7108)
         );
  AND4_X2 U7674 ( .A1(n8945), .A2(n8946), .A3(n8947), .A4(n8948), .ZN(n7110)
         );
  AND4_X2 U7675 ( .A1(n8913), .A2(n8914), .A3(n8915), .A4(n8916), .ZN(n7111)
         );
  AND4_X2 U7676 ( .A1(n8977), .A2(n8978), .A3(n8979), .A4(n8980), .ZN(n7112)
         );
  AND4_X2 U7677 ( .A1(n8881), .A2(n8882), .A3(n8883), .A4(n8884), .ZN(n7113)
         );
  AND4_X2 U7678 ( .A1(n9199), .A2(n9200), .A3(n9201), .A4(n9202), .ZN(n7114)
         );
  AND4_X2 U7679 ( .A1(n9103), .A2(n9104), .A3(n9105), .A4(n9106), .ZN(n7116)
         );
  AND4_X2 U7680 ( .A1(n7377), .A2(n7378), .A3(n7379), .A4(n7380), .ZN(n7119)
         );
  AND4_X2 U7681 ( .A1(n7505), .A2(n7506), .A3(n7507), .A4(n7508), .ZN(n7120)
         );
  AND4_X2 U7682 ( .A1(n8593), .A2(n8594), .A3(n8595), .A4(n8596), .ZN(n7121)
         );
  AND4_X2 U7683 ( .A1(n7729), .A2(n7730), .A3(n7731), .A4(n7732), .ZN(n7131)
         );
  AOI221_X2 U7684 ( .B1(pipeline_PC_DX[28]), .B2(n6958), .C1(
        pipeline_handler_PC[28]), .C2(n6630), .A(n12427), .ZN(n12428) );
  AND4_X2 U7685 ( .A1(n8529), .A2(n8530), .A3(n8531), .A4(n8532), .ZN(n7140)
         );
  AND4_X2 U7686 ( .A1(n8657), .A2(n8658), .A3(n8659), .A4(n8660), .ZN(n7142)
         );
  AND4_X2 U7687 ( .A1(n7441), .A2(n7442), .A3(n7443), .A4(n7444), .ZN(n7145)
         );
  AND4_X2 U7688 ( .A1(n8433), .A2(n8434), .A3(n8435), .A4(n8436), .ZN(n7147)
         );
  OAI22_X2 U7689 ( .A1(n9440), .A2(n6787), .B1(n12933), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[9]) );
  NOR2_X2 U7690 ( .A1(n7149), .A2(n7150), .ZN(n9141) );
  NOR2_X2 U7691 ( .A1(n7151), .A2(n7152), .ZN(n9013) );
  NOR2_X2 U7692 ( .A1(n7153), .A2(n7154), .ZN(n8951) );
  NOR2_X2 U7693 ( .A1(n7155), .A2(n7156), .ZN(n9077) );
  NOR2_X2 U7694 ( .A1(n7157), .A2(n7158), .ZN(n8631) );
  NOR2_X2 U7695 ( .A1(n7159), .A2(n7160), .ZN(n8695) );
  NOR2_X2 U7696 ( .A1(n7161), .A2(n7162), .ZN(n8791) );
  AOI21_X1 U7697 ( .B1(imem_hready), .B2(n12395), .A(pipeline_ctrl_replay_IF), 
        .ZN(n12406) );
  OAI21_X1 U7698 ( .B1(n636), .B2(n12557), .A(n12552), .ZN(
        pipeline_PCmux_offset[15]) );
  NAND2_X2 U7699 ( .A1(n9820), .A2(pipeline_imm_31_), .ZN(n9967) );
  OAI21_X1 U7700 ( .B1(n637), .B2(n12557), .A(n12552), .ZN(
        pipeline_PCmux_offset[16]) );
  OAI21_X1 U7701 ( .B1(imem_hready), .B2(n10094), .A(n10092), .ZN(n10385) );
  OAI21_X2 U7702 ( .B1(n800), .B2(n11179), .A(n10345), .ZN(n6049) );
  INV_X4 U7703 ( .A(n9465), .ZN(n9464) );
  INV_X4 U7704 ( .A(n11262), .ZN(n9465) );
  OR2_X1 U7705 ( .A1(n789), .A2(dmem_hready), .ZN(n9610) );
  AND3_X2 U7706 ( .A1(n7054), .A2(n8214), .A3(n6641), .ZN(n7166) );
  AND3_X2 U7707 ( .A1(n8223), .A2(n702), .A3(n8214), .ZN(n7167) );
  OR2_X1 U7708 ( .A1(ext_interrupts[16]), .A2(ext_interrupts[9]), .ZN(n9605)
         );
  OAI22_X2 U7709 ( .A1(n723), .A2(n9445), .B1(n12505), .B2(n9443), .ZN(
        pipeline_alu_src_a[8]) );
  NOR3_X2 U7710 ( .A1(pipeline_csr_N2405), .A2(n9629), .A3(pipeline_csr_N2407), 
        .ZN(n7177) );
  AND4_X2 U7711 ( .A1(n9647), .A2(n9646), .A3(n9645), .A4(n9644), .ZN(n7178)
         );
  AOI21_X2 U7712 ( .B1(htif_pcr_req_data[0]), .B2(n13131), .A(n11277), .ZN(
        n11278) );
  AOI21_X2 U7713 ( .B1(htif_pcr_req_data[2]), .B2(n13131), .A(n10414), .ZN(
        n10415) );
  AND4_X2 U7714 ( .A1(n9634), .A2(n6794), .A3(n10248), .A4(n7182), .ZN(n7180)
         );
  AND2_X1 U7715 ( .A1(n6711), .A2(n10336), .ZN(n7181) );
  AOI22_X2 U7716 ( .A1(pipeline_md_N24), .A2(n136), .B1(n135), .B2(n13145), 
        .ZN(n152) );
  AND2_X1 U7717 ( .A1(n6810), .A2(n9642), .ZN(n7183) );
  OR2_X1 U7718 ( .A1(n10188), .A2(n7184), .ZN(n10187) );
  INV_X4 U7719 ( .A(n12615), .ZN(n9491) );
  AND4_X2 U7720 ( .A1(n10687), .A2(n10686), .A3(n10685), .A4(n10684), .ZN(
        n7185) );
  NAND2_X2 U7721 ( .A1(pipeline_alu_out_WB[0]), .A2(n12936), .ZN(n12891) );
  AOI22_X2 U7722 ( .A1(n150), .A2(pipeline_md_N24), .B1(n149), .B2(n13145), 
        .ZN(n151) );
  NAND2_X2 U7723 ( .A1(n12850), .A2(n12940), .ZN(n12893) );
  NAND2_X2 U7724 ( .A1(pipeline_alu_out_WB[0]), .A2(pipeline_alu_out_WB[1]), 
        .ZN(n12981) );
  NAND2_X2 U7725 ( .A1(pipeline_alu_out_WB[1]), .A2(n12937), .ZN(n12979) );
  AND4_X2 U7726 ( .A1(n10738), .A2(n10737), .A3(n10736), .A4(n10735), .ZN(
        n7186) );
  AOI21_X2 U7727 ( .B1(n6748), .B2(n7051), .A(htif_reset), .ZN(n12600) );
  AND3_X2 U7728 ( .A1(n10904), .A2(n10903), .A3(n10902), .ZN(n7187) );
  AND3_X2 U7729 ( .A1(n11011), .A2(n11010), .A3(n11009), .ZN(n7188) );
  AND3_X2 U7730 ( .A1(n11121), .A2(n11120), .A3(n11119), .ZN(n7189) );
  AND2_X1 U7731 ( .A1(n10349), .A2(n13130), .ZN(n7190) );
  INV_X4 U7732 ( .A(n9533), .ZN(n9532) );
  INV_X4 U7733 ( .A(n2009), .ZN(n9533) );
  AND4_X2 U7734 ( .A1(n10958), .A2(n10957), .A3(n10956), .A4(n10955), .ZN(
        n7194) );
  AND4_X2 U7735 ( .A1(n11065), .A2(n11064), .A3(n11063), .A4(n11062), .ZN(
        n7195) );
  AND4_X2 U7736 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(
        n7196) );
  AND4_X2 U7737 ( .A1(n11150), .A2(n11149), .A3(n11148), .A4(n11147), .ZN(
        n7197) );
  AND4_X2 U7738 ( .A1(n11038), .A2(n11037), .A3(n11036), .A4(n11035), .ZN(
        n7198) );
  AND4_X2 U7739 ( .A1(n10877), .A2(n10876), .A3(n10875), .A4(n10874), .ZN(
        n7199) );
  AND4_X2 U7740 ( .A1(n10931), .A2(n10930), .A3(n10929), .A4(n10928), .ZN(
        n7200) );
  AND4_X2 U7741 ( .A1(n10985), .A2(n10984), .A3(n10983), .A4(n10982), .ZN(
        n7201) );
  AND4_X2 U7742 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n7202) );
  AND4_X2 U7743 ( .A1(n10850), .A2(n10849), .A3(n10848), .A4(n10847), .ZN(
        n7203) );
  AND4_X2 U7744 ( .A1(n10765), .A2(n10764), .A3(n10763), .A4(n10762), .ZN(
        n7204) );
  AND4_X2 U7745 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n7205) );
  AND4_X2 U7746 ( .A1(n10659), .A2(n10658), .A3(n10657), .A4(n10656), .ZN(
        n7206) );
  AND4_X2 U7747 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        n7207) );
  AND4_X2 U7748 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n7208) );
  AND4_X2 U7749 ( .A1(n10475), .A2(n10474), .A3(n10473), .A4(n10472), .ZN(
        n7209) );
  AND4_X2 U7750 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n7210) );
  AND4_X2 U7751 ( .A1(n10257), .A2(n10256), .A3(n10255), .A4(n10254), .ZN(
        n7211) );
  AND4_X2 U7752 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n7212) );
  AND3_X2 U7753 ( .A1(n10631), .A2(n10630), .A3(n10629), .ZN(n7213) );
  AND3_X2 U7754 ( .A1(n10299), .A2(n10298), .A3(n10297), .ZN(n7214) );
  NAND2_X2 U7755 ( .A1(n9535), .A2(pipeline_wb_src_sel_WB_0_), .ZN(n12985) );
  INV_X4 U7756 ( .A(htif_reset), .ZN(n13130) );
  INV_X4 U7757 ( .A(n9519), .ZN(n9518) );
  INV_X4 U7758 ( .A(n13029), .ZN(n9519) );
  AND2_X1 U7759 ( .A1(n12388), .A2(pipeline_ctrl_had_ex_WB), .ZN(n7215) );
  OAI222_X2 U7760 ( .A1(n503), .A2(n4229), .B1(n511), .B2(n4230), .C1(n13144), 
        .C2(n527), .ZN(dmem_hwdata[24]) );
  OAI222_X2 U7761 ( .A1(n504), .A2(n4229), .B1(n512), .B2(n4230), .C1(n13144), 
        .C2(n528), .ZN(dmem_hwdata[25]) );
  OAI222_X2 U7762 ( .A1(n505), .A2(n4229), .B1(n513), .B2(n4230), .C1(n13144), 
        .C2(n529), .ZN(dmem_hwdata[26]) );
  OAI222_X2 U7763 ( .A1(n506), .A2(n4229), .B1(n514), .B2(n4230), .C1(n13144), 
        .C2(n530), .ZN(dmem_hwdata[27]) );
  OAI222_X2 U7764 ( .A1(n507), .A2(n4229), .B1(n515), .B2(n4230), .C1(n13144), 
        .C2(n531), .ZN(dmem_hwdata[28]) );
  OAI222_X2 U7765 ( .A1(n508), .A2(n4229), .B1(n516), .B2(n4230), .C1(n13144), 
        .C2(n532), .ZN(dmem_hwdata[29]) );
  OAI222_X2 U7766 ( .A1(n509), .A2(n4229), .B1(n517), .B2(n4230), .C1(n13144), 
        .C2(n533), .ZN(dmem_hwdata[30]) );
  OAI222_X2 U7767 ( .A1(n510), .A2(n4229), .B1(n518), .B2(n4230), .C1(n13144), 
        .C2(n534), .ZN(dmem_hwdata[31]) );
  OR4_X1 U7768 ( .A1(pipeline_ctrl_prev_ex_code_WB[0]), .A2(
        pipeline_ctrl_prev_ex_code_WB[3]), .A3(n12292), .A4(n7216), .ZN(n11192) );
  OAI21_X2 U7769 ( .B1(htif_pcr_req_ready), .B2(n4205), .A(n4206), .ZN(n6368)
         );
  AOI221_X2 U7770 ( .B1(pipeline_regfile_data[928]), .B2(n6728), .C1(
        pipeline_regfile_data[672]), .C2(n6720), .A(n7221), .ZN(n7220) );
  OAI22_X2 U7771 ( .A1(n7222), .A2(n6695), .B1(n7223), .B2(n6663), .ZN(n7221)
         );
  AND2_X1 U7772 ( .A1(n7224), .A2(n7225), .ZN(n7223) );
  AOI221_X2 U7773 ( .B1(pipeline_regfile_data[352]), .B2(n8249), .C1(
        pipeline_regfile_data[288]), .C2(n8252), .A(n7227), .ZN(n7225) );
  NAND2_X2 U7774 ( .A1(n7228), .A2(n7229), .ZN(n7227) );
  NAND2_X2 U7775 ( .A1(pipeline_regfile_data[480]), .A2(n8254), .ZN(n7229) );
  NAND2_X2 U7776 ( .A1(pipeline_regfile_data[416]), .A2(n8257), .ZN(n7228) );
  AOI221_X2 U7777 ( .B1(pipeline_regfile_data[320]), .B2(n8261), .C1(
        pipeline_regfile_data[256]), .C2(n8263), .A(n7230), .ZN(n7224) );
  NAND2_X2 U7778 ( .A1(n7231), .A2(n7232), .ZN(n7230) );
  NAND2_X2 U7779 ( .A1(pipeline_regfile_data[448]), .A2(n8266), .ZN(n7232) );
  NAND2_X2 U7780 ( .A1(pipeline_regfile_data[384]), .A2(n8271), .ZN(n7231) );
  AND2_X1 U7781 ( .A1(n7233), .A2(n7234), .ZN(n7222) );
  AOI221_X2 U7782 ( .B1(pipeline_regfile_data[96]), .B2(n8249), .C1(
        pipeline_regfile_data[32]), .C2(n8253), .A(n7235), .ZN(n7234) );
  NAND2_X2 U7783 ( .A1(n7236), .A2(n7237), .ZN(n7235) );
  NAND2_X2 U7784 ( .A1(pipeline_regfile_data[224]), .A2(n8255), .ZN(n7237) );
  NAND2_X2 U7785 ( .A1(pipeline_regfile_data[160]), .A2(n8257), .ZN(n7236) );
  AOI221_X2 U7786 ( .B1(pipeline_regfile_data[64]), .B2(n8261), .C1(
        pipeline_regfile_data[0]), .C2(n8264), .A(n7238), .ZN(n7233) );
  NAND2_X2 U7787 ( .A1(n7239), .A2(n7240), .ZN(n7238) );
  NAND2_X2 U7788 ( .A1(pipeline_regfile_data[192]), .A2(n8266), .ZN(n7240) );
  NAND2_X2 U7789 ( .A1(pipeline_regfile_data[128]), .A2(n8269), .ZN(n7239) );
  AOI221_X2 U7790 ( .B1(pipeline_regfile_data[992]), .B2(n6725), .C1(
        pipeline_regfile_data[736]), .C2(n6721), .A(n7241), .ZN(n7219) );
  INV_X4 U7791 ( .A(n7242), .ZN(n7241) );
  AOI221_X2 U7792 ( .B1(pipeline_regfile_data[544]), .B2(n6726), .C1(
        pipeline_regfile_data[800]), .C2(n6722), .A(n7243), .ZN(n7242) );
  AND2_X1 U7793 ( .A1(pipeline_regfile_data[608]), .A2(n6730), .ZN(n7243) );
  NAND2_X2 U7794 ( .A1(n7245), .A2(n7246), .ZN(n7244) );
  NAND2_X2 U7795 ( .A1(pipeline_regfile_data[640]), .A2(n6731), .ZN(n7246) );
  NAND2_X2 U7796 ( .A1(pipeline_regfile_data[864]), .A2(n6732), .ZN(n7245) );
  AOI221_X2 U7797 ( .B1(pipeline_regfile_data[512]), .B2(n6719), .C1(
        pipeline_regfile_data[960]), .C2(n6723), .A(n7247), .ZN(n7217) );
  INV_X4 U7798 ( .A(n7248), .ZN(n7247) );
  AOI221_X2 U7799 ( .B1(pipeline_regfile_data[768]), .B2(n6727), .C1(
        pipeline_regfile_data[576]), .C2(n6724), .A(n7249), .ZN(n7248) );
  AND2_X1 U7800 ( .A1(pipeline_regfile_data[832]), .A2(n6729), .ZN(n7249) );
  AOI221_X2 U7801 ( .B1(pipeline_regfile_data[929]), .B2(n6728), .C1(
        pipeline_regfile_data[673]), .C2(n6720), .A(n7254), .ZN(n7253) );
  OAI22_X2 U7802 ( .A1(n7255), .A2(n6695), .B1(n7256), .B2(n6663), .ZN(n7254)
         );
  NAND2_X2 U7803 ( .A1(pipeline_regfile_data[481]), .A2(n8256), .ZN(n7260) );
  NAND2_X2 U7804 ( .A1(pipeline_regfile_data[417]), .A2(n8257), .ZN(n7259) );
  AOI221_X2 U7805 ( .B1(pipeline_regfile_data[321]), .B2(n8261), .C1(
        pipeline_regfile_data[257]), .C2(n8263), .A(n7261), .ZN(n7257) );
  NAND2_X2 U7806 ( .A1(n7262), .A2(n7263), .ZN(n7261) );
  NAND2_X2 U7807 ( .A1(pipeline_regfile_data[449]), .A2(n8266), .ZN(n7263) );
  NAND2_X2 U7808 ( .A1(pipeline_regfile_data[385]), .A2(n8271), .ZN(n7262) );
  AOI221_X2 U7809 ( .B1(pipeline_regfile_data[97]), .B2(n8249), .C1(
        pipeline_regfile_data[33]), .C2(n8252), .A(n7266), .ZN(n7265) );
  NAND2_X2 U7810 ( .A1(n7267), .A2(n7268), .ZN(n7266) );
  NAND2_X2 U7811 ( .A1(pipeline_regfile_data[225]), .A2(n8254), .ZN(n7268) );
  NAND2_X2 U7812 ( .A1(pipeline_regfile_data[161]), .A2(n8257), .ZN(n7267) );
  AOI221_X2 U7813 ( .B1(pipeline_regfile_data[65]), .B2(n8261), .C1(
        pipeline_regfile_data[1]), .C2(n8264), .A(n7269), .ZN(n7264) );
  NAND2_X2 U7814 ( .A1(n7270), .A2(n7271), .ZN(n7269) );
  NAND2_X2 U7815 ( .A1(pipeline_regfile_data[193]), .A2(n8266), .ZN(n7271) );
  NAND2_X2 U7816 ( .A1(pipeline_regfile_data[129]), .A2(n8271), .ZN(n7270) );
  AOI221_X2 U7817 ( .B1(pipeline_regfile_data[993]), .B2(n6725), .C1(
        pipeline_regfile_data[737]), .C2(n6721), .A(n7272), .ZN(n7252) );
  INV_X4 U7818 ( .A(n7273), .ZN(n7272) );
  AOI221_X2 U7819 ( .B1(pipeline_regfile_data[545]), .B2(n6726), .C1(
        pipeline_regfile_data[801]), .C2(n6722), .A(n7274), .ZN(n7273) );
  AND2_X1 U7820 ( .A1(pipeline_regfile_data[609]), .A2(n6730), .ZN(n7274) );
  AOI221_X2 U7821 ( .B1(pipeline_regfile_data[705]), .B2(n6734), .C1(
        pipeline_regfile_data[897]), .C2(n6733), .A(n7275), .ZN(n7251) );
  NAND2_X2 U7822 ( .A1(n7276), .A2(n7277), .ZN(n7275) );
  NAND2_X2 U7823 ( .A1(pipeline_regfile_data[641]), .A2(n6731), .ZN(n7277) );
  NAND2_X2 U7824 ( .A1(pipeline_regfile_data[865]), .A2(n6732), .ZN(n7276) );
  AOI221_X2 U7825 ( .B1(pipeline_regfile_data[513]), .B2(n6719), .C1(
        pipeline_regfile_data[961]), .C2(n6723), .A(n7278), .ZN(n7250) );
  INV_X4 U7826 ( .A(n7279), .ZN(n7278) );
  AOI221_X2 U7827 ( .B1(pipeline_regfile_data[769]), .B2(n6727), .C1(
        pipeline_regfile_data[577]), .C2(n6724), .A(n7280), .ZN(n7279) );
  AND2_X1 U7828 ( .A1(pipeline_regfile_data[833]), .A2(n6729), .ZN(n7280) );
  AOI221_X2 U7829 ( .B1(pipeline_regfile_data[930]), .B2(n6728), .C1(
        pipeline_regfile_data[674]), .C2(n6720), .A(n7285), .ZN(n7284) );
  OAI22_X2 U7830 ( .A1(n7286), .A2(n6695), .B1(n7287), .B2(n6663), .ZN(n7285)
         );
  AND2_X1 U7831 ( .A1(n7288), .A2(n7289), .ZN(n7287) );
  AOI221_X2 U7832 ( .B1(pipeline_regfile_data[354]), .B2(n8249), .C1(
        pipeline_regfile_data[290]), .C2(n8253), .A(n7290), .ZN(n7289) );
  NAND2_X2 U7833 ( .A1(n7291), .A2(n7292), .ZN(n7290) );
  NAND2_X2 U7834 ( .A1(pipeline_regfile_data[482]), .A2(n8255), .ZN(n7292) );
  NAND2_X2 U7835 ( .A1(pipeline_regfile_data[418]), .A2(n8257), .ZN(n7291) );
  AOI221_X2 U7836 ( .B1(pipeline_regfile_data[322]), .B2(n8261), .C1(
        pipeline_regfile_data[258]), .C2(n8264), .A(n7293), .ZN(n7288) );
  NAND2_X2 U7837 ( .A1(n7294), .A2(n7295), .ZN(n7293) );
  NAND2_X2 U7838 ( .A1(pipeline_regfile_data[450]), .A2(n8266), .ZN(n7295) );
  NAND2_X2 U7839 ( .A1(pipeline_regfile_data[386]), .A2(n8269), .ZN(n7294) );
  AND2_X1 U7840 ( .A1(n7296), .A2(n7297), .ZN(n7286) );
  AOI221_X2 U7841 ( .B1(pipeline_regfile_data[98]), .B2(n8249), .C1(
        pipeline_regfile_data[34]), .C2(n8253), .A(n7298), .ZN(n7297) );
  NAND2_X2 U7842 ( .A1(n7299), .A2(n7300), .ZN(n7298) );
  NAND2_X2 U7843 ( .A1(pipeline_regfile_data[226]), .A2(n8255), .ZN(n7300) );
  NAND2_X2 U7844 ( .A1(pipeline_regfile_data[162]), .A2(n8257), .ZN(n7299) );
  AOI221_X2 U7845 ( .B1(pipeline_regfile_data[66]), .B2(n8261), .C1(
        pipeline_regfile_data[2]), .C2(n8264), .A(n7301), .ZN(n7296) );
  NAND2_X2 U7846 ( .A1(n7302), .A2(n7303), .ZN(n7301) );
  NAND2_X2 U7847 ( .A1(pipeline_regfile_data[194]), .A2(n8266), .ZN(n7303) );
  NAND2_X2 U7848 ( .A1(pipeline_regfile_data[130]), .A2(n8269), .ZN(n7302) );
  AOI221_X2 U7849 ( .B1(pipeline_regfile_data[994]), .B2(n6725), .C1(
        pipeline_regfile_data[738]), .C2(n6721), .A(n7304), .ZN(n7283) );
  INV_X4 U7850 ( .A(n7305), .ZN(n7304) );
  AOI221_X2 U7851 ( .B1(pipeline_regfile_data[546]), .B2(n6726), .C1(
        pipeline_regfile_data[802]), .C2(n6722), .A(n7306), .ZN(n7305) );
  AND2_X1 U7852 ( .A1(pipeline_regfile_data[610]), .A2(n6730), .ZN(n7306) );
  NAND2_X2 U7853 ( .A1(n7308), .A2(n7309), .ZN(n7307) );
  NAND2_X2 U7854 ( .A1(pipeline_regfile_data[642]), .A2(n6731), .ZN(n7309) );
  NAND2_X2 U7855 ( .A1(pipeline_regfile_data[866]), .A2(n6732), .ZN(n7308) );
  AOI221_X2 U7856 ( .B1(pipeline_regfile_data[514]), .B2(n6719), .C1(
        pipeline_regfile_data[962]), .C2(n6723), .A(n7310), .ZN(n7281) );
  INV_X4 U7857 ( .A(n7311), .ZN(n7310) );
  AOI221_X2 U7858 ( .B1(pipeline_regfile_data[770]), .B2(n6727), .C1(
        pipeline_regfile_data[578]), .C2(n6724), .A(n7312), .ZN(n7311) );
  AND2_X1 U7859 ( .A1(pipeline_regfile_data[834]), .A2(n6729), .ZN(n7312) );
  AOI221_X2 U7860 ( .B1(pipeline_regfile_data[931]), .B2(n6728), .C1(
        pipeline_regfile_data[675]), .C2(n6720), .A(n7317), .ZN(n7316) );
  OAI22_X2 U7861 ( .A1(n7318), .A2(n6695), .B1(n7319), .B2(n6663), .ZN(n7317)
         );
  AND2_X1 U7862 ( .A1(n7320), .A2(n7321), .ZN(n7319) );
  NAND2_X2 U7863 ( .A1(n7323), .A2(n7324), .ZN(n7322) );
  NAND2_X2 U7864 ( .A1(pipeline_regfile_data[483]), .A2(n8255), .ZN(n7324) );
  NAND2_X2 U7865 ( .A1(pipeline_regfile_data[419]), .A2(n8257), .ZN(n7323) );
  AOI221_X2 U7866 ( .B1(pipeline_regfile_data[323]), .B2(n8261), .C1(
        pipeline_regfile_data[259]), .C2(n8262), .A(n7325), .ZN(n7320) );
  NAND2_X2 U7867 ( .A1(n7326), .A2(n7327), .ZN(n7325) );
  NAND2_X2 U7868 ( .A1(pipeline_regfile_data[451]), .A2(n8266), .ZN(n7327) );
  NAND2_X2 U7869 ( .A1(pipeline_regfile_data[387]), .A2(n8271), .ZN(n7326) );
  AND2_X1 U7870 ( .A1(n7328), .A2(n7329), .ZN(n7318) );
  AOI221_X2 U7871 ( .B1(pipeline_regfile_data[99]), .B2(n8249), .C1(
        pipeline_regfile_data[35]), .C2(n8253), .A(n7330), .ZN(n7329) );
  NAND2_X2 U7872 ( .A1(n7331), .A2(n7332), .ZN(n7330) );
  NAND2_X2 U7873 ( .A1(pipeline_regfile_data[227]), .A2(n8255), .ZN(n7332) );
  NAND2_X2 U7874 ( .A1(pipeline_regfile_data[163]), .A2(n8257), .ZN(n7331) );
  AOI221_X2 U7875 ( .B1(pipeline_regfile_data[67]), .B2(n8261), .C1(
        pipeline_regfile_data[3]), .C2(n8263), .A(n7333), .ZN(n7328) );
  NAND2_X2 U7876 ( .A1(n7334), .A2(n7335), .ZN(n7333) );
  NAND2_X2 U7877 ( .A1(pipeline_regfile_data[195]), .A2(n8266), .ZN(n7335) );
  NAND2_X2 U7878 ( .A1(pipeline_regfile_data[131]), .A2(n8270), .ZN(n7334) );
  AOI221_X2 U7879 ( .B1(pipeline_regfile_data[995]), .B2(n6725), .C1(
        pipeline_regfile_data[739]), .C2(n6721), .A(n7336), .ZN(n7315) );
  INV_X4 U7880 ( .A(n7337), .ZN(n7336) );
  AOI221_X2 U7881 ( .B1(pipeline_regfile_data[547]), .B2(n6726), .C1(
        pipeline_regfile_data[803]), .C2(n6722), .A(n7338), .ZN(n7337) );
  AND2_X1 U7882 ( .A1(pipeline_regfile_data[611]), .A2(n6730), .ZN(n7338) );
  AOI221_X2 U7883 ( .B1(pipeline_regfile_data[707]), .B2(n6734), .C1(
        pipeline_regfile_data[899]), .C2(n6733), .A(n7339), .ZN(n7314) );
  NAND2_X2 U7884 ( .A1(n7340), .A2(n7341), .ZN(n7339) );
  NAND2_X2 U7885 ( .A1(pipeline_regfile_data[643]), .A2(n6731), .ZN(n7341) );
  NAND2_X2 U7886 ( .A1(pipeline_regfile_data[867]), .A2(n6732), .ZN(n7340) );
  AOI221_X2 U7887 ( .B1(pipeline_regfile_data[515]), .B2(n6719), .C1(
        pipeline_regfile_data[963]), .C2(n6723), .A(n7342), .ZN(n7313) );
  INV_X4 U7888 ( .A(n7343), .ZN(n7342) );
  AOI221_X2 U7889 ( .B1(pipeline_regfile_data[771]), .B2(n6727), .C1(
        pipeline_regfile_data[579]), .C2(n6724), .A(n7344), .ZN(n7343) );
  AND2_X1 U7890 ( .A1(pipeline_regfile_data[835]), .A2(n6729), .ZN(n7344) );
  AOI221_X2 U7891 ( .B1(pipeline_regfile_data[932]), .B2(n6728), .C1(
        pipeline_regfile_data[676]), .C2(n6720), .A(n7349), .ZN(n7348) );
  OAI22_X2 U7892 ( .A1(n7350), .A2(n6695), .B1(n7351), .B2(n6663), .ZN(n7349)
         );
  AOI221_X2 U7893 ( .B1(pipeline_regfile_data[356]), .B2(n8249), .C1(
        pipeline_regfile_data[292]), .C2(n8253), .A(n7354), .ZN(n7353) );
  NAND2_X2 U7894 ( .A1(n7355), .A2(n7356), .ZN(n7354) );
  NAND2_X2 U7895 ( .A1(pipeline_regfile_data[484]), .A2(n8256), .ZN(n7356) );
  NAND2_X2 U7896 ( .A1(pipeline_regfile_data[420]), .A2(n8257), .ZN(n7355) );
  AOI221_X2 U7897 ( .B1(pipeline_regfile_data[324]), .B2(n8261), .C1(
        pipeline_regfile_data[260]), .C2(n8262), .A(n7357), .ZN(n7352) );
  NAND2_X2 U7898 ( .A1(n7358), .A2(n7359), .ZN(n7357) );
  NAND2_X2 U7899 ( .A1(pipeline_regfile_data[452]), .A2(n8266), .ZN(n7359) );
  NAND2_X2 U7900 ( .A1(pipeline_regfile_data[388]), .A2(n8271), .ZN(n7358) );
  AND2_X1 U7901 ( .A1(n7360), .A2(n7361), .ZN(n7350) );
  AOI221_X2 U7902 ( .B1(pipeline_regfile_data[100]), .B2(n8249), .C1(
        pipeline_regfile_data[36]), .C2(n8252), .A(n7362), .ZN(n7361) );
  NAND2_X2 U7903 ( .A1(n7363), .A2(n7364), .ZN(n7362) );
  NAND2_X2 U7904 ( .A1(pipeline_regfile_data[228]), .A2(n8255), .ZN(n7364) );
  NAND2_X2 U7905 ( .A1(pipeline_regfile_data[164]), .A2(n8257), .ZN(n7363) );
  AOI221_X2 U7906 ( .B1(pipeline_regfile_data[68]), .B2(n8261), .C1(
        pipeline_regfile_data[4]), .C2(n8265), .A(n7365), .ZN(n7360) );
  NAND2_X2 U7907 ( .A1(n7366), .A2(n7367), .ZN(n7365) );
  NAND2_X2 U7908 ( .A1(pipeline_regfile_data[196]), .A2(n8266), .ZN(n7367) );
  NAND2_X2 U7909 ( .A1(pipeline_regfile_data[132]), .A2(n8271), .ZN(n7366) );
  AOI221_X2 U7910 ( .B1(pipeline_regfile_data[996]), .B2(n6725), .C1(
        pipeline_regfile_data[740]), .C2(n6721), .A(n7368), .ZN(n7347) );
  INV_X4 U7911 ( .A(n7369), .ZN(n7368) );
  AOI221_X2 U7912 ( .B1(pipeline_regfile_data[548]), .B2(n6726), .C1(
        pipeline_regfile_data[804]), .C2(n6722), .A(n7370), .ZN(n7369) );
  AND2_X1 U7913 ( .A1(pipeline_regfile_data[612]), .A2(n6730), .ZN(n7370) );
  AOI221_X2 U7914 ( .B1(pipeline_regfile_data[708]), .B2(n6734), .C1(
        pipeline_regfile_data[900]), .C2(n6733), .A(n7371), .ZN(n7346) );
  NAND2_X2 U7915 ( .A1(n7372), .A2(n7373), .ZN(n7371) );
  NAND2_X2 U7916 ( .A1(pipeline_regfile_data[644]), .A2(n6731), .ZN(n7373) );
  NAND2_X2 U7917 ( .A1(pipeline_regfile_data[868]), .A2(n6732), .ZN(n7372) );
  AOI221_X2 U7918 ( .B1(pipeline_regfile_data[516]), .B2(n6719), .C1(
        pipeline_regfile_data[964]), .C2(n6723), .A(n7374), .ZN(n7345) );
  AOI221_X2 U7919 ( .B1(pipeline_regfile_data[772]), .B2(n6727), .C1(
        pipeline_regfile_data[580]), .C2(n6724), .A(n7376), .ZN(n7375) );
  AOI221_X2 U7920 ( .B1(pipeline_regfile_data[933]), .B2(n6728), .C1(
        pipeline_regfile_data[677]), .C2(n6720), .A(n7381), .ZN(n7380) );
  OAI22_X2 U7921 ( .A1(n7382), .A2(n6695), .B1(n7383), .B2(n6663), .ZN(n7381)
         );
  AND2_X1 U7922 ( .A1(n7384), .A2(n7385), .ZN(n7383) );
  NAND2_X2 U7923 ( .A1(n7387), .A2(n7388), .ZN(n7386) );
  NAND2_X2 U7924 ( .A1(pipeline_regfile_data[485]), .A2(n8255), .ZN(n7388) );
  NAND2_X2 U7925 ( .A1(pipeline_regfile_data[421]), .A2(n8257), .ZN(n7387) );
  AOI221_X2 U7926 ( .B1(pipeline_regfile_data[325]), .B2(n8261), .C1(
        pipeline_regfile_data[261]), .C2(n8265), .A(n7389), .ZN(n7384) );
  NAND2_X2 U7927 ( .A1(n7390), .A2(n7391), .ZN(n7389) );
  NAND2_X2 U7928 ( .A1(pipeline_regfile_data[453]), .A2(n8266), .ZN(n7391) );
  NAND2_X2 U7929 ( .A1(pipeline_regfile_data[389]), .A2(n8270), .ZN(n7390) );
  AND2_X1 U7930 ( .A1(n7392), .A2(n7393), .ZN(n7382) );
  NAND2_X2 U7931 ( .A1(n7395), .A2(n7396), .ZN(n7394) );
  NAND2_X2 U7932 ( .A1(pipeline_regfile_data[229]), .A2(n8255), .ZN(n7396) );
  NAND2_X2 U7933 ( .A1(pipeline_regfile_data[165]), .A2(n8257), .ZN(n7395) );
  AOI221_X2 U7934 ( .B1(pipeline_regfile_data[69]), .B2(n8261), .C1(
        pipeline_regfile_data[5]), .C2(n8265), .A(n7397), .ZN(n7392) );
  NAND2_X2 U7935 ( .A1(n7398), .A2(n7399), .ZN(n7397) );
  NAND2_X2 U7936 ( .A1(pipeline_regfile_data[197]), .A2(n8266), .ZN(n7399) );
  NAND2_X2 U7937 ( .A1(pipeline_regfile_data[133]), .A2(n8269), .ZN(n7398) );
  AOI221_X2 U7938 ( .B1(pipeline_regfile_data[997]), .B2(n6725), .C1(
        pipeline_regfile_data[741]), .C2(n6721), .A(n7400), .ZN(n7379) );
  INV_X4 U7939 ( .A(n7401), .ZN(n7400) );
  AOI221_X2 U7940 ( .B1(pipeline_regfile_data[549]), .B2(n6726), .C1(
        pipeline_regfile_data[805]), .C2(n6722), .A(n7402), .ZN(n7401) );
  AND2_X1 U7941 ( .A1(pipeline_regfile_data[613]), .A2(n6730), .ZN(n7402) );
  NAND2_X2 U7942 ( .A1(n7404), .A2(n7405), .ZN(n7403) );
  NAND2_X2 U7943 ( .A1(pipeline_regfile_data[645]), .A2(n6731), .ZN(n7405) );
  NAND2_X2 U7944 ( .A1(pipeline_regfile_data[869]), .A2(n6732), .ZN(n7404) );
  AOI221_X2 U7945 ( .B1(pipeline_regfile_data[517]), .B2(n6719), .C1(
        pipeline_regfile_data[965]), .C2(n6723), .A(n7406), .ZN(n7377) );
  INV_X4 U7946 ( .A(n7407), .ZN(n7406) );
  AOI221_X2 U7947 ( .B1(pipeline_regfile_data[773]), .B2(n6727), .C1(
        pipeline_regfile_data[581]), .C2(n6724), .A(n7408), .ZN(n7407) );
  AND2_X1 U7948 ( .A1(pipeline_regfile_data[837]), .A2(n6729), .ZN(n7408) );
  AOI221_X2 U7949 ( .B1(pipeline_regfile_data[934]), .B2(n6728), .C1(
        pipeline_regfile_data[678]), .C2(n6720), .A(n7413), .ZN(n7412) );
  OAI22_X2 U7950 ( .A1(n7414), .A2(n6695), .B1(n7415), .B2(n6663), .ZN(n7413)
         );
  AND2_X1 U7951 ( .A1(n7416), .A2(n7417), .ZN(n7415) );
  AOI221_X2 U7952 ( .B1(pipeline_regfile_data[358]), .B2(n8249), .C1(
        pipeline_regfile_data[294]), .C2(n8253), .A(n7418), .ZN(n7417) );
  NAND2_X2 U7953 ( .A1(n7419), .A2(n7420), .ZN(n7418) );
  NAND2_X2 U7954 ( .A1(pipeline_regfile_data[486]), .A2(n8255), .ZN(n7420) );
  NAND2_X2 U7955 ( .A1(pipeline_regfile_data[422]), .A2(n8257), .ZN(n7419) );
  AOI221_X2 U7956 ( .B1(pipeline_regfile_data[326]), .B2(n8261), .C1(
        pipeline_regfile_data[262]), .C2(n8263), .A(n7421), .ZN(n7416) );
  NAND2_X2 U7957 ( .A1(n7422), .A2(n7423), .ZN(n7421) );
  NAND2_X2 U7958 ( .A1(pipeline_regfile_data[454]), .A2(n8266), .ZN(n7423) );
  NAND2_X2 U7959 ( .A1(pipeline_regfile_data[390]), .A2(n8269), .ZN(n7422) );
  AND2_X1 U7960 ( .A1(n7424), .A2(n7425), .ZN(n7414) );
  AOI221_X2 U7961 ( .B1(pipeline_regfile_data[102]), .B2(n8248), .C1(
        pipeline_regfile_data[38]), .C2(n8253), .A(n7426), .ZN(n7425) );
  NAND2_X2 U7962 ( .A1(n7427), .A2(n7428), .ZN(n7426) );
  NAND2_X2 U7963 ( .A1(pipeline_regfile_data[230]), .A2(n8255), .ZN(n7428) );
  NAND2_X2 U7964 ( .A1(pipeline_regfile_data[166]), .A2(n8257), .ZN(n7427) );
  AOI221_X2 U7965 ( .B1(pipeline_regfile_data[70]), .B2(n8260), .C1(
        pipeline_regfile_data[6]), .C2(n8263), .A(n7429), .ZN(n7424) );
  NAND2_X2 U7966 ( .A1(n7430), .A2(n7431), .ZN(n7429) );
  NAND2_X2 U7967 ( .A1(pipeline_regfile_data[198]), .A2(n8266), .ZN(n7431) );
  NAND2_X2 U7968 ( .A1(pipeline_regfile_data[134]), .A2(n8271), .ZN(n7430) );
  AOI221_X2 U7969 ( .B1(pipeline_regfile_data[998]), .B2(n6725), .C1(
        pipeline_regfile_data[742]), .C2(n6721), .A(n7432), .ZN(n7411) );
  INV_X4 U7970 ( .A(n7433), .ZN(n7432) );
  AOI221_X2 U7971 ( .B1(pipeline_regfile_data[550]), .B2(n6726), .C1(
        pipeline_regfile_data[806]), .C2(n6722), .A(n7434), .ZN(n7433) );
  AND2_X1 U7972 ( .A1(pipeline_regfile_data[614]), .A2(n6730), .ZN(n7434) );
  NAND2_X2 U7973 ( .A1(n7436), .A2(n7437), .ZN(n7435) );
  NAND2_X2 U7974 ( .A1(pipeline_regfile_data[646]), .A2(n6731), .ZN(n7437) );
  NAND2_X2 U7975 ( .A1(pipeline_regfile_data[870]), .A2(n6732), .ZN(n7436) );
  AOI221_X2 U7976 ( .B1(pipeline_regfile_data[518]), .B2(n6719), .C1(
        pipeline_regfile_data[966]), .C2(n6723), .A(n7438), .ZN(n7409) );
  INV_X4 U7977 ( .A(n7439), .ZN(n7438) );
  AOI221_X2 U7978 ( .B1(pipeline_regfile_data[774]), .B2(n6727), .C1(
        pipeline_regfile_data[582]), .C2(n6724), .A(n7440), .ZN(n7439) );
  AND2_X1 U7979 ( .A1(pipeline_regfile_data[838]), .A2(n6729), .ZN(n7440) );
  AOI221_X2 U7980 ( .B1(pipeline_regfile_data[935]), .B2(n6728), .C1(
        pipeline_regfile_data[679]), .C2(n6720), .A(n7445), .ZN(n7444) );
  OAI22_X2 U7981 ( .A1(n7446), .A2(n6695), .B1(n7447), .B2(n6663), .ZN(n7445)
         );
  AND2_X1 U7982 ( .A1(n7448), .A2(n7449), .ZN(n7447) );
  AOI221_X2 U7983 ( .B1(pipeline_regfile_data[359]), .B2(n8248), .C1(
        pipeline_regfile_data[295]), .C2(n8253), .A(n7450), .ZN(n7449) );
  NAND2_X2 U7984 ( .A1(n7451), .A2(n7452), .ZN(n7450) );
  NAND2_X2 U7985 ( .A1(pipeline_regfile_data[423]), .A2(n8257), .ZN(n7451) );
  AOI221_X2 U7986 ( .B1(pipeline_regfile_data[327]), .B2(n8260), .C1(
        pipeline_regfile_data[263]), .C2(n8265), .A(n7453), .ZN(n7448) );
  NAND2_X2 U7987 ( .A1(n7454), .A2(n7455), .ZN(n7453) );
  NAND2_X2 U7988 ( .A1(pipeline_regfile_data[455]), .A2(n8268), .ZN(n7455) );
  NAND2_X2 U7989 ( .A1(pipeline_regfile_data[391]), .A2(n8270), .ZN(n7454) );
  AND2_X1 U7990 ( .A1(n7456), .A2(n7457), .ZN(n7446) );
  NAND2_X2 U7991 ( .A1(n7459), .A2(n7460), .ZN(n7458) );
  NAND2_X2 U7992 ( .A1(pipeline_regfile_data[231]), .A2(n8254), .ZN(n7460) );
  NAND2_X2 U7993 ( .A1(pipeline_regfile_data[167]), .A2(n8257), .ZN(n7459) );
  AOI221_X2 U7994 ( .B1(pipeline_regfile_data[71]), .B2(n8260), .C1(
        pipeline_regfile_data[7]), .C2(n8264), .A(n7461), .ZN(n7456) );
  NAND2_X2 U7995 ( .A1(n7462), .A2(n7463), .ZN(n7461) );
  NAND2_X2 U7996 ( .A1(pipeline_regfile_data[199]), .A2(n8268), .ZN(n7463) );
  NAND2_X2 U7997 ( .A1(pipeline_regfile_data[135]), .A2(n8270), .ZN(n7462) );
  AOI221_X2 U7998 ( .B1(pipeline_regfile_data[999]), .B2(n6725), .C1(
        pipeline_regfile_data[743]), .C2(n6721), .A(n7464), .ZN(n7443) );
  INV_X4 U7999 ( .A(n7465), .ZN(n7464) );
  AOI221_X2 U8000 ( .B1(pipeline_regfile_data[551]), .B2(n6726), .C1(
        pipeline_regfile_data[807]), .C2(n6722), .A(n7466), .ZN(n7465) );
  AND2_X1 U8001 ( .A1(pipeline_regfile_data[615]), .A2(n6730), .ZN(n7466) );
  NAND2_X2 U8002 ( .A1(n7468), .A2(n7469), .ZN(n7467) );
  NAND2_X2 U8003 ( .A1(pipeline_regfile_data[647]), .A2(n6731), .ZN(n7469) );
  NAND2_X2 U8004 ( .A1(pipeline_regfile_data[871]), .A2(n6732), .ZN(n7468) );
  AOI221_X2 U8005 ( .B1(pipeline_regfile_data[519]), .B2(n6719), .C1(
        pipeline_regfile_data[967]), .C2(n6723), .A(n7470), .ZN(n7441) );
  INV_X4 U8006 ( .A(n7471), .ZN(n7470) );
  AOI221_X2 U8007 ( .B1(pipeline_regfile_data[775]), .B2(n6727), .C1(
        pipeline_regfile_data[583]), .C2(n6724), .A(n7472), .ZN(n7471) );
  AND2_X1 U8008 ( .A1(pipeline_regfile_data[839]), .A2(n6729), .ZN(n7472) );
  AOI221_X2 U8009 ( .B1(pipeline_regfile_data[936]), .B2(n6728), .C1(
        pipeline_regfile_data[680]), .C2(n6720), .A(n7477), .ZN(n7476) );
  OAI22_X2 U8010 ( .A1(n7478), .A2(n6695), .B1(n7479), .B2(n6663), .ZN(n7477)
         );
  NAND2_X2 U8011 ( .A1(n7483), .A2(n7484), .ZN(n7482) );
  NAND2_X2 U8012 ( .A1(pipeline_regfile_data[488]), .A2(n8254), .ZN(n7484) );
  NAND2_X2 U8013 ( .A1(pipeline_regfile_data[424]), .A2(n8257), .ZN(n7483) );
  AOI221_X2 U8014 ( .B1(pipeline_regfile_data[328]), .B2(n8260), .C1(
        pipeline_regfile_data[264]), .C2(n8263), .A(n7485), .ZN(n7480) );
  NAND2_X2 U8015 ( .A1(n7486), .A2(n7487), .ZN(n7485) );
  NAND2_X2 U8016 ( .A1(pipeline_regfile_data[456]), .A2(n8268), .ZN(n7487) );
  NAND2_X2 U8017 ( .A1(pipeline_regfile_data[392]), .A2(n8269), .ZN(n7486) );
  AND2_X1 U8018 ( .A1(n7488), .A2(n7489), .ZN(n7478) );
  NAND2_X2 U8019 ( .A1(n7491), .A2(n7492), .ZN(n7490) );
  NAND2_X2 U8020 ( .A1(pipeline_regfile_data[232]), .A2(n8254), .ZN(n7492) );
  NAND2_X2 U8021 ( .A1(pipeline_regfile_data[168]), .A2(n8257), .ZN(n7491) );
  AOI221_X2 U8022 ( .B1(pipeline_regfile_data[72]), .B2(n8260), .C1(
        pipeline_regfile_data[8]), .C2(n8265), .A(n7493), .ZN(n7488) );
  NAND2_X2 U8023 ( .A1(n7494), .A2(n7495), .ZN(n7493) );
  NAND2_X2 U8024 ( .A1(pipeline_regfile_data[200]), .A2(n8268), .ZN(n7495) );
  NAND2_X2 U8025 ( .A1(pipeline_regfile_data[136]), .A2(n8269), .ZN(n7494) );
  AOI221_X2 U8026 ( .B1(pipeline_regfile_data[1000]), .B2(n6725), .C1(
        pipeline_regfile_data[744]), .C2(n6721), .A(n7496), .ZN(n7475) );
  INV_X4 U8027 ( .A(n7497), .ZN(n7496) );
  AOI221_X2 U8028 ( .B1(pipeline_regfile_data[552]), .B2(n6726), .C1(
        pipeline_regfile_data[808]), .C2(n6722), .A(n7498), .ZN(n7497) );
  AND2_X1 U8029 ( .A1(pipeline_regfile_data[616]), .A2(n6730), .ZN(n7498) );
  NAND2_X2 U8030 ( .A1(n7500), .A2(n7501), .ZN(n7499) );
  NAND2_X2 U8031 ( .A1(pipeline_regfile_data[648]), .A2(n6731), .ZN(n7501) );
  NAND2_X2 U8032 ( .A1(pipeline_regfile_data[872]), .A2(n6732), .ZN(n7500) );
  AOI221_X2 U8033 ( .B1(pipeline_regfile_data[520]), .B2(n6719), .C1(
        pipeline_regfile_data[968]), .C2(n6723), .A(n7502), .ZN(n7473) );
  INV_X4 U8034 ( .A(n7503), .ZN(n7502) );
  AOI221_X2 U8035 ( .B1(pipeline_regfile_data[776]), .B2(n6727), .C1(
        pipeline_regfile_data[584]), .C2(n6724), .A(n7504), .ZN(n7503) );
  AND2_X1 U8036 ( .A1(pipeline_regfile_data[840]), .A2(n6729), .ZN(n7504) );
  AOI221_X2 U8037 ( .B1(pipeline_regfile_data[937]), .B2(n6728), .C1(
        pipeline_regfile_data[681]), .C2(n6720), .A(n7509), .ZN(n7508) );
  OAI22_X2 U8038 ( .A1(n7510), .A2(n6695), .B1(n7511), .B2(n6663), .ZN(n7509)
         );
  AND2_X1 U8039 ( .A1(n7512), .A2(n7513), .ZN(n7511) );
  NAND2_X2 U8040 ( .A1(n7515), .A2(n7516), .ZN(n7514) );
  NAND2_X2 U8041 ( .A1(pipeline_regfile_data[489]), .A2(n8254), .ZN(n7516) );
  NAND2_X2 U8042 ( .A1(pipeline_regfile_data[425]), .A2(n8257), .ZN(n7515) );
  AOI221_X2 U8043 ( .B1(pipeline_regfile_data[329]), .B2(n8260), .C1(
        pipeline_regfile_data[265]), .C2(n8265), .A(n7517), .ZN(n7512) );
  NAND2_X2 U8044 ( .A1(n7518), .A2(n7519), .ZN(n7517) );
  NAND2_X2 U8045 ( .A1(pipeline_regfile_data[457]), .A2(n8266), .ZN(n7519) );
  NAND2_X2 U8046 ( .A1(pipeline_regfile_data[393]), .A2(n8270), .ZN(n7518) );
  AND2_X1 U8047 ( .A1(n7520), .A2(n7521), .ZN(n7510) );
  NAND2_X2 U8048 ( .A1(n7523), .A2(n7524), .ZN(n7522) );
  NAND2_X2 U8049 ( .A1(pipeline_regfile_data[233]), .A2(n8254), .ZN(n7524) );
  NAND2_X2 U8050 ( .A1(pipeline_regfile_data[169]), .A2(n8257), .ZN(n7523) );
  AOI221_X2 U8051 ( .B1(pipeline_regfile_data[73]), .B2(n8260), .C1(
        pipeline_regfile_data[9]), .C2(n8264), .A(n7525), .ZN(n7520) );
  NAND2_X2 U8052 ( .A1(n7526), .A2(n7527), .ZN(n7525) );
  NAND2_X2 U8053 ( .A1(pipeline_regfile_data[201]), .A2(n8268), .ZN(n7527) );
  NAND2_X2 U8054 ( .A1(pipeline_regfile_data[137]), .A2(n8270), .ZN(n7526) );
  AOI221_X2 U8055 ( .B1(pipeline_regfile_data[1001]), .B2(n6725), .C1(
        pipeline_regfile_data[745]), .C2(n6721), .A(n7528), .ZN(n7507) );
  INV_X4 U8056 ( .A(n7529), .ZN(n7528) );
  AOI221_X2 U8057 ( .B1(pipeline_regfile_data[553]), .B2(n6726), .C1(
        pipeline_regfile_data[809]), .C2(n6722), .A(n7530), .ZN(n7529) );
  AND2_X1 U8058 ( .A1(pipeline_regfile_data[617]), .A2(n6730), .ZN(n7530) );
  NAND2_X2 U8059 ( .A1(n7532), .A2(n7533), .ZN(n7531) );
  NAND2_X2 U8060 ( .A1(pipeline_regfile_data[649]), .A2(n6731), .ZN(n7533) );
  NAND2_X2 U8061 ( .A1(pipeline_regfile_data[873]), .A2(n6732), .ZN(n7532) );
  AOI221_X2 U8062 ( .B1(pipeline_regfile_data[521]), .B2(n6719), .C1(
        pipeline_regfile_data[969]), .C2(n6723), .A(n7534), .ZN(n7505) );
  INV_X4 U8063 ( .A(n7535), .ZN(n7534) );
  AOI221_X2 U8064 ( .B1(pipeline_regfile_data[777]), .B2(n6727), .C1(
        pipeline_regfile_data[585]), .C2(n6724), .A(n7536), .ZN(n7535) );
  AND2_X1 U8065 ( .A1(pipeline_regfile_data[841]), .A2(n6729), .ZN(n7536) );
  AOI221_X2 U8066 ( .B1(pipeline_regfile_data[938]), .B2(n6728), .C1(
        pipeline_regfile_data[682]), .C2(n6720), .A(n7541), .ZN(n7540) );
  OAI22_X2 U8067 ( .A1(n7542), .A2(n6695), .B1(n7543), .B2(n6663), .ZN(n7541)
         );
  AND2_X1 U8068 ( .A1(n7544), .A2(n7545), .ZN(n7543) );
  AOI221_X2 U8069 ( .B1(pipeline_regfile_data[362]), .B2(n8248), .C1(
        pipeline_regfile_data[298]), .C2(n8253), .A(n7546), .ZN(n7545) );
  NAND2_X2 U8070 ( .A1(n7547), .A2(n7548), .ZN(n7546) );
  NAND2_X2 U8071 ( .A1(pipeline_regfile_data[426]), .A2(n8257), .ZN(n7547) );
  AOI221_X2 U8072 ( .B1(pipeline_regfile_data[330]), .B2(n8260), .C1(
        pipeline_regfile_data[266]), .C2(n8263), .A(n7549), .ZN(n7544) );
  NAND2_X2 U8073 ( .A1(n7550), .A2(n7551), .ZN(n7549) );
  NAND2_X2 U8074 ( .A1(pipeline_regfile_data[458]), .A2(n8268), .ZN(n7551) );
  NAND2_X2 U8075 ( .A1(pipeline_regfile_data[394]), .A2(n8270), .ZN(n7550) );
  AND2_X1 U8076 ( .A1(n7552), .A2(n7553), .ZN(n7542) );
  NAND2_X2 U8077 ( .A1(n7555), .A2(n7556), .ZN(n7554) );
  NAND2_X2 U8078 ( .A1(pipeline_regfile_data[234]), .A2(n8254), .ZN(n7556) );
  NAND2_X2 U8079 ( .A1(pipeline_regfile_data[170]), .A2(n8257), .ZN(n7555) );
  AOI221_X2 U8080 ( .B1(pipeline_regfile_data[74]), .B2(n8260), .C1(
        pipeline_regfile_data[10]), .C2(n8264), .A(n7557), .ZN(n7552) );
  NAND2_X2 U8081 ( .A1(n7558), .A2(n7559), .ZN(n7557) );
  NAND2_X2 U8082 ( .A1(pipeline_regfile_data[202]), .A2(n8268), .ZN(n7559) );
  NAND2_X2 U8083 ( .A1(pipeline_regfile_data[138]), .A2(n8271), .ZN(n7558) );
  AOI221_X2 U8084 ( .B1(pipeline_regfile_data[1002]), .B2(n6725), .C1(
        pipeline_regfile_data[746]), .C2(n6721), .A(n7560), .ZN(n7539) );
  INV_X4 U8085 ( .A(n7561), .ZN(n7560) );
  AOI221_X2 U8086 ( .B1(pipeline_regfile_data[554]), .B2(n6726), .C1(
        pipeline_regfile_data[810]), .C2(n6722), .A(n7562), .ZN(n7561) );
  AND2_X1 U8087 ( .A1(pipeline_regfile_data[618]), .A2(n6730), .ZN(n7562) );
  NAND2_X2 U8088 ( .A1(n7564), .A2(n7565), .ZN(n7563) );
  NAND2_X2 U8089 ( .A1(pipeline_regfile_data[650]), .A2(n6731), .ZN(n7565) );
  NAND2_X2 U8090 ( .A1(pipeline_regfile_data[874]), .A2(n6732), .ZN(n7564) );
  AOI221_X2 U8091 ( .B1(pipeline_regfile_data[522]), .B2(n6719), .C1(
        pipeline_regfile_data[970]), .C2(n6723), .A(n7566), .ZN(n7537) );
  INV_X4 U8092 ( .A(n7567), .ZN(n7566) );
  AOI221_X2 U8093 ( .B1(pipeline_regfile_data[778]), .B2(n6727), .C1(
        pipeline_regfile_data[586]), .C2(n6724), .A(n7568), .ZN(n7567) );
  AND2_X1 U8094 ( .A1(pipeline_regfile_data[842]), .A2(n6729), .ZN(n7568) );
  AOI221_X2 U8095 ( .B1(pipeline_regfile_data[939]), .B2(n6728), .C1(
        pipeline_regfile_data[683]), .C2(n6720), .A(n7573), .ZN(n7572) );
  OAI22_X2 U8096 ( .A1(n7574), .A2(n6695), .B1(n7575), .B2(n6663), .ZN(n7573)
         );
  AND2_X1 U8097 ( .A1(n7576), .A2(n7577), .ZN(n7575) );
  AOI221_X2 U8098 ( .B1(pipeline_regfile_data[363]), .B2(n8248), .C1(
        pipeline_regfile_data[299]), .C2(n8253), .A(n7578), .ZN(n7577) );
  NAND2_X2 U8099 ( .A1(n7579), .A2(n7580), .ZN(n7578) );
  NAND2_X2 U8100 ( .A1(pipeline_regfile_data[491]), .A2(n8254), .ZN(n7580) );
  NAND2_X2 U8101 ( .A1(pipeline_regfile_data[427]), .A2(n8257), .ZN(n7579) );
  AOI221_X2 U8102 ( .B1(pipeline_regfile_data[331]), .B2(n8260), .C1(
        pipeline_regfile_data[267]), .C2(n8265), .A(n7581), .ZN(n7576) );
  NAND2_X2 U8103 ( .A1(n7582), .A2(n7583), .ZN(n7581) );
  NAND2_X2 U8104 ( .A1(pipeline_regfile_data[459]), .A2(n8268), .ZN(n7583) );
  NAND2_X2 U8105 ( .A1(pipeline_regfile_data[395]), .A2(n8269), .ZN(n7582) );
  AND2_X1 U8106 ( .A1(n7584), .A2(n7585), .ZN(n7574) );
  NAND2_X2 U8107 ( .A1(n7587), .A2(n7588), .ZN(n7586) );
  NAND2_X2 U8108 ( .A1(pipeline_regfile_data[235]), .A2(n8254), .ZN(n7588) );
  NAND2_X2 U8109 ( .A1(pipeline_regfile_data[171]), .A2(n8257), .ZN(n7587) );
  AOI221_X2 U8110 ( .B1(pipeline_regfile_data[75]), .B2(n8260), .C1(
        pipeline_regfile_data[11]), .C2(n8264), .A(n7589), .ZN(n7584) );
  NAND2_X2 U8111 ( .A1(n7590), .A2(n7591), .ZN(n7589) );
  NAND2_X2 U8112 ( .A1(pipeline_regfile_data[203]), .A2(n8266), .ZN(n7591) );
  NAND2_X2 U8113 ( .A1(pipeline_regfile_data[139]), .A2(n8271), .ZN(n7590) );
  AOI221_X2 U8114 ( .B1(pipeline_regfile_data[1003]), .B2(n6725), .C1(
        pipeline_regfile_data[747]), .C2(n6721), .A(n7592), .ZN(n7571) );
  INV_X4 U8115 ( .A(n7593), .ZN(n7592) );
  AOI221_X2 U8116 ( .B1(pipeline_regfile_data[555]), .B2(n6726), .C1(
        pipeline_regfile_data[811]), .C2(n6722), .A(n7594), .ZN(n7593) );
  AND2_X1 U8117 ( .A1(pipeline_regfile_data[619]), .A2(n6730), .ZN(n7594) );
  NAND2_X2 U8118 ( .A1(n7596), .A2(n7597), .ZN(n7595) );
  NAND2_X2 U8119 ( .A1(pipeline_regfile_data[651]), .A2(n6731), .ZN(n7597) );
  NAND2_X2 U8120 ( .A1(pipeline_regfile_data[875]), .A2(n6732), .ZN(n7596) );
  AOI221_X2 U8121 ( .B1(pipeline_regfile_data[523]), .B2(n6719), .C1(
        pipeline_regfile_data[971]), .C2(n6723), .A(n7598), .ZN(n7569) );
  INV_X4 U8122 ( .A(n7599), .ZN(n7598) );
  AOI221_X2 U8123 ( .B1(pipeline_regfile_data[779]), .B2(n6727), .C1(
        pipeline_regfile_data[587]), .C2(n6724), .A(n7600), .ZN(n7599) );
  AND2_X1 U8124 ( .A1(pipeline_regfile_data[843]), .A2(n6729), .ZN(n7600) );
  AOI221_X2 U8125 ( .B1(pipeline_regfile_data[940]), .B2(n6728), .C1(
        pipeline_regfile_data[684]), .C2(n6720), .A(n7605), .ZN(n7604) );
  OAI22_X2 U8126 ( .A1(n7606), .A2(n6695), .B1(n7607), .B2(n6663), .ZN(n7605)
         );
  AOI221_X2 U8127 ( .B1(pipeline_regfile_data[364]), .B2(n8248), .C1(
        pipeline_regfile_data[300]), .C2(n8252), .A(n7610), .ZN(n7609) );
  NAND2_X2 U8128 ( .A1(n7611), .A2(n7612), .ZN(n7610) );
  NAND2_X2 U8129 ( .A1(pipeline_regfile_data[492]), .A2(n8254), .ZN(n7612) );
  NAND2_X2 U8130 ( .A1(pipeline_regfile_data[428]), .A2(n8257), .ZN(n7611) );
  AOI221_X2 U8131 ( .B1(pipeline_regfile_data[332]), .B2(n8260), .C1(
        pipeline_regfile_data[268]), .C2(n8263), .A(n7613), .ZN(n7608) );
  NAND2_X2 U8132 ( .A1(n7614), .A2(n7615), .ZN(n7613) );
  NAND2_X2 U8133 ( .A1(pipeline_regfile_data[460]), .A2(n8268), .ZN(n7615) );
  NAND2_X2 U8134 ( .A1(pipeline_regfile_data[396]), .A2(n8271), .ZN(n7614) );
  AND2_X1 U8135 ( .A1(n7616), .A2(n7617), .ZN(n7606) );
  AOI221_X2 U8136 ( .B1(pipeline_regfile_data[108]), .B2(n8248), .C1(
        pipeline_regfile_data[44]), .C2(n8252), .A(n7618), .ZN(n7617) );
  NAND2_X2 U8137 ( .A1(n7619), .A2(n7620), .ZN(n7618) );
  NAND2_X2 U8138 ( .A1(pipeline_regfile_data[236]), .A2(n8254), .ZN(n7620) );
  NAND2_X2 U8139 ( .A1(pipeline_regfile_data[172]), .A2(n8257), .ZN(n7619) );
  AOI221_X2 U8140 ( .B1(pipeline_regfile_data[76]), .B2(n8260), .C1(
        pipeline_regfile_data[12]), .C2(n8265), .A(n7621), .ZN(n7616) );
  NAND2_X2 U8141 ( .A1(n7622), .A2(n7623), .ZN(n7621) );
  NAND2_X2 U8142 ( .A1(pipeline_regfile_data[204]), .A2(n8268), .ZN(n7623) );
  NAND2_X2 U8143 ( .A1(pipeline_regfile_data[140]), .A2(n8271), .ZN(n7622) );
  AOI221_X2 U8144 ( .B1(pipeline_regfile_data[1004]), .B2(n6725), .C1(
        pipeline_regfile_data[748]), .C2(n6721), .A(n7624), .ZN(n7603) );
  INV_X4 U8145 ( .A(n7625), .ZN(n7624) );
  AOI221_X2 U8146 ( .B1(pipeline_regfile_data[556]), .B2(n6726), .C1(
        pipeline_regfile_data[812]), .C2(n6722), .A(n7626), .ZN(n7625) );
  AND2_X1 U8147 ( .A1(pipeline_regfile_data[620]), .A2(n6730), .ZN(n7626) );
  AOI221_X2 U8148 ( .B1(pipeline_regfile_data[716]), .B2(n6734), .C1(
        pipeline_regfile_data[908]), .C2(n6733), .A(n7627), .ZN(n7602) );
  NAND2_X2 U8149 ( .A1(n7628), .A2(n7629), .ZN(n7627) );
  NAND2_X2 U8150 ( .A1(pipeline_regfile_data[652]), .A2(n6731), .ZN(n7629) );
  NAND2_X2 U8151 ( .A1(pipeline_regfile_data[876]), .A2(n6732), .ZN(n7628) );
  AOI221_X2 U8152 ( .B1(pipeline_regfile_data[524]), .B2(n6719), .C1(
        pipeline_regfile_data[972]), .C2(n6723), .A(n7630), .ZN(n7601) );
  INV_X4 U8153 ( .A(n7631), .ZN(n7630) );
  AOI221_X2 U8154 ( .B1(pipeline_regfile_data[780]), .B2(n6727), .C1(
        pipeline_regfile_data[588]), .C2(n6724), .A(n7632), .ZN(n7631) );
  AND2_X1 U8155 ( .A1(pipeline_regfile_data[844]), .A2(n6729), .ZN(n7632) );
  AOI221_X2 U8156 ( .B1(pipeline_regfile_data[941]), .B2(n6728), .C1(
        pipeline_regfile_data[685]), .C2(n6720), .A(n7637), .ZN(n7636) );
  OAI22_X2 U8157 ( .A1(n7638), .A2(n6695), .B1(n7639), .B2(n6663), .ZN(n7637)
         );
  AND2_X1 U8158 ( .A1(n7640), .A2(n7641), .ZN(n7639) );
  AOI221_X2 U8159 ( .B1(pipeline_regfile_data[365]), .B2(n8247), .C1(
        pipeline_regfile_data[301]), .C2(n8253), .A(n7642), .ZN(n7641) );
  NAND2_X2 U8160 ( .A1(n7643), .A2(n7644), .ZN(n7642) );
  NAND2_X2 U8161 ( .A1(pipeline_regfile_data[493]), .A2(n8254), .ZN(n7644) );
  NAND2_X2 U8162 ( .A1(pipeline_regfile_data[429]), .A2(n8257), .ZN(n7643) );
  AOI221_X2 U8163 ( .B1(pipeline_regfile_data[333]), .B2(n8259), .C1(
        pipeline_regfile_data[269]), .C2(n8265), .A(n7645), .ZN(n7640) );
  NAND2_X2 U8164 ( .A1(n7646), .A2(n7647), .ZN(n7645) );
  NAND2_X2 U8165 ( .A1(pipeline_regfile_data[461]), .A2(n8266), .ZN(n7647) );
  NAND2_X2 U8166 ( .A1(pipeline_regfile_data[397]), .A2(n8269), .ZN(n7646) );
  AND2_X1 U8167 ( .A1(n7648), .A2(n7649), .ZN(n7638) );
  AOI221_X2 U8168 ( .B1(pipeline_regfile_data[109]), .B2(n8247), .C1(
        pipeline_regfile_data[45]), .C2(n8252), .A(n7650), .ZN(n7649) );
  NAND2_X2 U8169 ( .A1(n7651), .A2(n7652), .ZN(n7650) );
  NAND2_X2 U8170 ( .A1(pipeline_regfile_data[237]), .A2(n8255), .ZN(n7652) );
  NAND2_X2 U8171 ( .A1(pipeline_regfile_data[173]), .A2(n8257), .ZN(n7651) );
  AOI221_X2 U8172 ( .B1(pipeline_regfile_data[77]), .B2(n8259), .C1(
        pipeline_regfile_data[13]), .C2(n8265), .A(n7653), .ZN(n7648) );
  NAND2_X2 U8173 ( .A1(n7654), .A2(n7655), .ZN(n7653) );
  NAND2_X2 U8174 ( .A1(pipeline_regfile_data[205]), .A2(n6599), .ZN(n7655) );
  NAND2_X2 U8175 ( .A1(pipeline_regfile_data[141]), .A2(n8269), .ZN(n7654) );
  AOI221_X2 U8176 ( .B1(pipeline_regfile_data[1005]), .B2(n6725), .C1(
        pipeline_regfile_data[749]), .C2(n6721), .A(n7656), .ZN(n7635) );
  INV_X4 U8177 ( .A(n7657), .ZN(n7656) );
  AOI221_X2 U8178 ( .B1(pipeline_regfile_data[557]), .B2(n6726), .C1(
        pipeline_regfile_data[813]), .C2(n6722), .A(n7658), .ZN(n7657) );
  AND2_X1 U8179 ( .A1(pipeline_regfile_data[621]), .A2(n6730), .ZN(n7658) );
  NAND2_X2 U8180 ( .A1(n7660), .A2(n7661), .ZN(n7659) );
  NAND2_X2 U8181 ( .A1(pipeline_regfile_data[653]), .A2(n6731), .ZN(n7661) );
  NAND2_X2 U8182 ( .A1(pipeline_regfile_data[877]), .A2(n6732), .ZN(n7660) );
  AOI221_X2 U8183 ( .B1(pipeline_regfile_data[525]), .B2(n6719), .C1(
        pipeline_regfile_data[973]), .C2(n6723), .A(n7662), .ZN(n7633) );
  INV_X4 U8184 ( .A(n7663), .ZN(n7662) );
  AOI221_X2 U8185 ( .B1(pipeline_regfile_data[781]), .B2(n6727), .C1(
        pipeline_regfile_data[589]), .C2(n6724), .A(n7664), .ZN(n7663) );
  AND2_X1 U8186 ( .A1(pipeline_regfile_data[845]), .A2(n6729), .ZN(n7664) );
  OAI22_X2 U8187 ( .A1(n7670), .A2(n6695), .B1(n7671), .B2(n6663), .ZN(n7669)
         );
  NAND2_X2 U8188 ( .A1(n7675), .A2(n7676), .ZN(n7674) );
  NAND2_X2 U8189 ( .A1(pipeline_regfile_data[494]), .A2(n8255), .ZN(n7676) );
  NAND2_X2 U8190 ( .A1(pipeline_regfile_data[430]), .A2(n8257), .ZN(n7675) );
  AOI221_X2 U8191 ( .B1(pipeline_regfile_data[334]), .B2(n8259), .C1(
        pipeline_regfile_data[270]), .C2(n8265), .A(n7677), .ZN(n7672) );
  NAND2_X2 U8192 ( .A1(n7678), .A2(n7679), .ZN(n7677) );
  NAND2_X2 U8193 ( .A1(pipeline_regfile_data[462]), .A2(n6599), .ZN(n7679) );
  NAND2_X2 U8194 ( .A1(pipeline_regfile_data[398]), .A2(n8269), .ZN(n7678) );
  AND2_X1 U8195 ( .A1(n7680), .A2(n7681), .ZN(n7670) );
  AOI221_X2 U8196 ( .B1(pipeline_regfile_data[110]), .B2(n8247), .C1(
        pipeline_regfile_data[46]), .C2(n8252), .A(n7682), .ZN(n7681) );
  NAND2_X2 U8197 ( .A1(n7683), .A2(n7684), .ZN(n7682) );
  NAND2_X2 U8198 ( .A1(pipeline_regfile_data[238]), .A2(n8255), .ZN(n7684) );
  NAND2_X2 U8199 ( .A1(pipeline_regfile_data[174]), .A2(n8257), .ZN(n7683) );
  AOI221_X2 U8200 ( .B1(pipeline_regfile_data[78]), .B2(n8259), .C1(
        pipeline_regfile_data[14]), .C2(n8263), .A(n7685), .ZN(n7680) );
  NAND2_X2 U8201 ( .A1(n7686), .A2(n7687), .ZN(n7685) );
  NAND2_X2 U8202 ( .A1(pipeline_regfile_data[206]), .A2(n6599), .ZN(n7687) );
  NAND2_X2 U8203 ( .A1(pipeline_regfile_data[142]), .A2(n8270), .ZN(n7686) );
  AOI221_X2 U8204 ( .B1(pipeline_regfile_data[1006]), .B2(n6725), .C1(
        pipeline_regfile_data[750]), .C2(n6721), .A(n7688), .ZN(n7667) );
  INV_X4 U8205 ( .A(n7689), .ZN(n7688) );
  AOI221_X2 U8206 ( .B1(pipeline_regfile_data[558]), .B2(n6726), .C1(
        pipeline_regfile_data[814]), .C2(n6722), .A(n7690), .ZN(n7689) );
  AND2_X1 U8207 ( .A1(pipeline_regfile_data[622]), .A2(n6730), .ZN(n7690) );
  NAND2_X2 U8208 ( .A1(n7692), .A2(n7693), .ZN(n7691) );
  NAND2_X2 U8209 ( .A1(pipeline_regfile_data[654]), .A2(n6731), .ZN(n7693) );
  NAND2_X2 U8210 ( .A1(pipeline_regfile_data[878]), .A2(n6732), .ZN(n7692) );
  AOI221_X2 U8211 ( .B1(pipeline_regfile_data[526]), .B2(n6719), .C1(
        pipeline_regfile_data[974]), .C2(n6723), .A(n7694), .ZN(n7665) );
  INV_X4 U8212 ( .A(n7695), .ZN(n7694) );
  AOI221_X2 U8213 ( .B1(pipeline_regfile_data[782]), .B2(n6727), .C1(
        pipeline_regfile_data[590]), .C2(n6724), .A(n7696), .ZN(n7695) );
  AND2_X1 U8214 ( .A1(pipeline_regfile_data[846]), .A2(n6729), .ZN(n7696) );
  AOI221_X2 U8215 ( .B1(pipeline_regfile_data[943]), .B2(n6728), .C1(
        pipeline_regfile_data[687]), .C2(n6720), .A(n7701), .ZN(n7700) );
  OAI22_X2 U8216 ( .A1(n7702), .A2(n6695), .B1(n7703), .B2(n6663), .ZN(n7701)
         );
  AND2_X1 U8217 ( .A1(n7704), .A2(n7705), .ZN(n7703) );
  AOI221_X2 U8218 ( .B1(pipeline_regfile_data[367]), .B2(n8247), .C1(
        pipeline_regfile_data[303]), .C2(n8253), .A(n7706), .ZN(n7705) );
  NAND2_X2 U8219 ( .A1(n7707), .A2(n7708), .ZN(n7706) );
  NAND2_X2 U8220 ( .A1(pipeline_regfile_data[495]), .A2(n8255), .ZN(n7708) );
  NAND2_X2 U8221 ( .A1(pipeline_regfile_data[431]), .A2(n8257), .ZN(n7707) );
  AOI221_X2 U8222 ( .B1(pipeline_regfile_data[335]), .B2(n8259), .C1(
        pipeline_regfile_data[271]), .C2(n8263), .A(n7709), .ZN(n7704) );
  NAND2_X2 U8223 ( .A1(n7710), .A2(n7711), .ZN(n7709) );
  NAND2_X2 U8224 ( .A1(pipeline_regfile_data[463]), .A2(n6599), .ZN(n7711) );
  NAND2_X2 U8225 ( .A1(pipeline_regfile_data[399]), .A2(n8269), .ZN(n7710) );
  AND2_X1 U8226 ( .A1(n7712), .A2(n7713), .ZN(n7702) );
  NAND2_X2 U8227 ( .A1(n7715), .A2(n7716), .ZN(n7714) );
  NAND2_X2 U8228 ( .A1(pipeline_regfile_data[239]), .A2(n8255), .ZN(n7716) );
  NAND2_X2 U8229 ( .A1(pipeline_regfile_data[175]), .A2(n8257), .ZN(n7715) );
  AOI221_X2 U8230 ( .B1(pipeline_regfile_data[79]), .B2(n8259), .C1(
        pipeline_regfile_data[15]), .C2(n8265), .A(n7717), .ZN(n7712) );
  NAND2_X2 U8231 ( .A1(n7718), .A2(n7719), .ZN(n7717) );
  NAND2_X2 U8232 ( .A1(pipeline_regfile_data[207]), .A2(n6599), .ZN(n7719) );
  NAND2_X2 U8233 ( .A1(pipeline_regfile_data[143]), .A2(n8271), .ZN(n7718) );
  AOI221_X2 U8234 ( .B1(pipeline_regfile_data[1007]), .B2(n6725), .C1(
        pipeline_regfile_data[751]), .C2(n6721), .A(n7720), .ZN(n7699) );
  INV_X4 U8235 ( .A(n7721), .ZN(n7720) );
  AOI221_X2 U8236 ( .B1(pipeline_regfile_data[559]), .B2(n6726), .C1(
        pipeline_regfile_data[815]), .C2(n6722), .A(n7722), .ZN(n7721) );
  AND2_X1 U8237 ( .A1(pipeline_regfile_data[623]), .A2(n6730), .ZN(n7722) );
  NAND2_X2 U8238 ( .A1(n7724), .A2(n7725), .ZN(n7723) );
  NAND2_X2 U8239 ( .A1(pipeline_regfile_data[655]), .A2(n6731), .ZN(n7725) );
  NAND2_X2 U8240 ( .A1(pipeline_regfile_data[879]), .A2(n6732), .ZN(n7724) );
  AOI221_X2 U8241 ( .B1(pipeline_regfile_data[527]), .B2(n6719), .C1(
        pipeline_regfile_data[975]), .C2(n6723), .A(n7726), .ZN(n7697) );
  INV_X4 U8242 ( .A(n7727), .ZN(n7726) );
  AOI221_X2 U8243 ( .B1(pipeline_regfile_data[783]), .B2(n6727), .C1(
        pipeline_regfile_data[591]), .C2(n6724), .A(n7728), .ZN(n7727) );
  AND2_X1 U8244 ( .A1(pipeline_regfile_data[847]), .A2(n6729), .ZN(n7728) );
  AOI221_X2 U8245 ( .B1(pipeline_regfile_data[944]), .B2(n6728), .C1(
        pipeline_regfile_data[688]), .C2(n6720), .A(n7733), .ZN(n7732) );
  OAI22_X2 U8246 ( .A1(n7734), .A2(n6695), .B1(n7735), .B2(n6663), .ZN(n7733)
         );
  AND2_X1 U8247 ( .A1(n7736), .A2(n7737), .ZN(n7735) );
  AOI221_X2 U8248 ( .B1(pipeline_regfile_data[368]), .B2(n8247), .C1(
        pipeline_regfile_data[304]), .C2(n8253), .A(n7738), .ZN(n7737) );
  NAND2_X2 U8249 ( .A1(n7739), .A2(n7740), .ZN(n7738) );
  NAND2_X2 U8250 ( .A1(pipeline_regfile_data[496]), .A2(n8255), .ZN(n7740) );
  NAND2_X2 U8251 ( .A1(pipeline_regfile_data[432]), .A2(n8257), .ZN(n7739) );
  AOI221_X2 U8252 ( .B1(pipeline_regfile_data[336]), .B2(n8259), .C1(
        pipeline_regfile_data[272]), .C2(n8263), .A(n7741), .ZN(n7736) );
  NAND2_X2 U8253 ( .A1(n7742), .A2(n7743), .ZN(n7741) );
  NAND2_X2 U8254 ( .A1(pipeline_regfile_data[464]), .A2(n6599), .ZN(n7743) );
  NAND2_X2 U8255 ( .A1(pipeline_regfile_data[400]), .A2(n8269), .ZN(n7742) );
  AND2_X1 U8256 ( .A1(n7744), .A2(n7745), .ZN(n7734) );
  AOI221_X2 U8257 ( .B1(pipeline_regfile_data[112]), .B2(n8247), .C1(
        pipeline_regfile_data[48]), .C2(n8253), .A(n7746), .ZN(n7745) );
  NAND2_X2 U8258 ( .A1(n7747), .A2(n7748), .ZN(n7746) );
  NAND2_X2 U8259 ( .A1(pipeline_regfile_data[240]), .A2(n8255), .ZN(n7748) );
  NAND2_X2 U8260 ( .A1(pipeline_regfile_data[176]), .A2(n8257), .ZN(n7747) );
  AOI221_X2 U8261 ( .B1(pipeline_regfile_data[80]), .B2(n8259), .C1(
        pipeline_regfile_data[16]), .C2(n8265), .A(n7749), .ZN(n7744) );
  NAND2_X2 U8262 ( .A1(n7750), .A2(n7751), .ZN(n7749) );
  NAND2_X2 U8263 ( .A1(pipeline_regfile_data[208]), .A2(n6599), .ZN(n7751) );
  NAND2_X2 U8264 ( .A1(pipeline_regfile_data[144]), .A2(n8269), .ZN(n7750) );
  AOI221_X2 U8265 ( .B1(pipeline_regfile_data[1008]), .B2(n6725), .C1(
        pipeline_regfile_data[752]), .C2(n6721), .A(n7752), .ZN(n7731) );
  INV_X4 U8266 ( .A(n7753), .ZN(n7752) );
  AOI221_X2 U8267 ( .B1(pipeline_regfile_data[560]), .B2(n6726), .C1(
        pipeline_regfile_data[816]), .C2(n6722), .A(n7754), .ZN(n7753) );
  AND2_X1 U8268 ( .A1(pipeline_regfile_data[624]), .A2(n6730), .ZN(n7754) );
  NAND2_X2 U8269 ( .A1(n7756), .A2(n7757), .ZN(n7755) );
  NAND2_X2 U8270 ( .A1(pipeline_regfile_data[656]), .A2(n6731), .ZN(n7757) );
  NAND2_X2 U8271 ( .A1(pipeline_regfile_data[880]), .A2(n6732), .ZN(n7756) );
  AOI221_X2 U8272 ( .B1(pipeline_regfile_data[528]), .B2(n6719), .C1(
        pipeline_regfile_data[976]), .C2(n6723), .A(n7758), .ZN(n7729) );
  INV_X4 U8273 ( .A(n7759), .ZN(n7758) );
  AOI221_X2 U8274 ( .B1(pipeline_regfile_data[784]), .B2(n6727), .C1(
        pipeline_regfile_data[592]), .C2(n6724), .A(n7760), .ZN(n7759) );
  AND2_X1 U8275 ( .A1(pipeline_regfile_data[848]), .A2(n6729), .ZN(n7760) );
  OAI22_X2 U8276 ( .A1(n7765), .A2(n6695), .B1(n7766), .B2(n6663), .ZN(n7764)
         );
  AND2_X1 U8277 ( .A1(n7767), .A2(n7768), .ZN(n7766) );
  NAND2_X2 U8278 ( .A1(n7770), .A2(n7771), .ZN(n7769) );
  NAND2_X2 U8279 ( .A1(pipeline_regfile_data[497]), .A2(n8255), .ZN(n7771) );
  NAND2_X2 U8280 ( .A1(pipeline_regfile_data[433]), .A2(n8257), .ZN(n7770) );
  AOI221_X2 U8281 ( .B1(pipeline_regfile_data[337]), .B2(n8259), .C1(
        pipeline_regfile_data[273]), .C2(n8263), .A(n7772), .ZN(n7767) );
  NAND2_X2 U8282 ( .A1(n7773), .A2(n7774), .ZN(n7772) );
  NAND2_X2 U8283 ( .A1(pipeline_regfile_data[465]), .A2(n6599), .ZN(n7774) );
  NAND2_X2 U8284 ( .A1(pipeline_regfile_data[401]), .A2(n8271), .ZN(n7773) );
  AND2_X1 U8285 ( .A1(n7775), .A2(n7776), .ZN(n7765) );
  NAND2_X2 U8286 ( .A1(n7778), .A2(n7779), .ZN(n7777) );
  NAND2_X2 U8287 ( .A1(pipeline_regfile_data[241]), .A2(n8255), .ZN(n7779) );
  NAND2_X2 U8288 ( .A1(pipeline_regfile_data[177]), .A2(n8257), .ZN(n7778) );
  AOI221_X2 U8289 ( .B1(pipeline_regfile_data[81]), .B2(n8259), .C1(
        pipeline_regfile_data[17]), .C2(n8262), .A(n7780), .ZN(n7775) );
  NAND2_X2 U8290 ( .A1(n7781), .A2(n7782), .ZN(n7780) );
  NAND2_X2 U8291 ( .A1(pipeline_regfile_data[209]), .A2(n6599), .ZN(n7782) );
  NAND2_X2 U8292 ( .A1(pipeline_regfile_data[145]), .A2(n8271), .ZN(n7781) );
  AOI221_X2 U8293 ( .B1(pipeline_regfile_data[1009]), .B2(n6725), .C1(
        pipeline_regfile_data[753]), .C2(n6721), .A(n7783), .ZN(n7763) );
  INV_X4 U8294 ( .A(n7784), .ZN(n7783) );
  AOI221_X2 U8295 ( .B1(pipeline_regfile_data[561]), .B2(n6726), .C1(
        pipeline_regfile_data[817]), .C2(n6722), .A(n7785), .ZN(n7784) );
  AND2_X1 U8296 ( .A1(pipeline_regfile_data[625]), .A2(n6730), .ZN(n7785) );
  AOI221_X2 U8297 ( .B1(pipeline_regfile_data[721]), .B2(n6734), .C1(
        pipeline_regfile_data[913]), .C2(n6733), .A(n7786), .ZN(n7762) );
  NAND2_X2 U8298 ( .A1(n7787), .A2(n7788), .ZN(n7786) );
  NAND2_X2 U8299 ( .A1(pipeline_regfile_data[657]), .A2(n6731), .ZN(n7788) );
  NAND2_X2 U8300 ( .A1(pipeline_regfile_data[881]), .A2(n6732), .ZN(n7787) );
  AOI221_X2 U8301 ( .B1(pipeline_regfile_data[529]), .B2(n6719), .C1(
        pipeline_regfile_data[977]), .C2(n6723), .A(n7789), .ZN(n7761) );
  INV_X4 U8302 ( .A(n7790), .ZN(n7789) );
  AOI221_X2 U8303 ( .B1(pipeline_regfile_data[785]), .B2(n6727), .C1(
        pipeline_regfile_data[593]), .C2(n6724), .A(n7791), .ZN(n7790) );
  AND2_X1 U8304 ( .A1(pipeline_regfile_data[849]), .A2(n6729), .ZN(n7791) );
  AOI221_X2 U8305 ( .B1(pipeline_regfile_data[946]), .B2(n6728), .C1(
        pipeline_regfile_data[690]), .C2(n6720), .A(n7796), .ZN(n7795) );
  OAI22_X2 U8306 ( .A1(n7797), .A2(n6695), .B1(n7798), .B2(n6663), .ZN(n7796)
         );
  AND2_X1 U8307 ( .A1(n7799), .A2(n7800), .ZN(n7798) );
  AOI221_X2 U8308 ( .B1(pipeline_regfile_data[370]), .B2(n8247), .C1(
        pipeline_regfile_data[306]), .C2(n8253), .A(n7801), .ZN(n7800) );
  NAND2_X2 U8309 ( .A1(n7802), .A2(n7803), .ZN(n7801) );
  NAND2_X2 U8310 ( .A1(pipeline_regfile_data[498]), .A2(n8255), .ZN(n7803) );
  NAND2_X2 U8311 ( .A1(pipeline_regfile_data[434]), .A2(n8257), .ZN(n7802) );
  AOI221_X2 U8312 ( .B1(pipeline_regfile_data[338]), .B2(n8259), .C1(
        pipeline_regfile_data[274]), .C2(n8263), .A(n7804), .ZN(n7799) );
  NAND2_X2 U8313 ( .A1(n7805), .A2(n7806), .ZN(n7804) );
  NAND2_X2 U8314 ( .A1(pipeline_regfile_data[466]), .A2(n6599), .ZN(n7806) );
  NAND2_X2 U8315 ( .A1(pipeline_regfile_data[402]), .A2(n8269), .ZN(n7805) );
  AND2_X1 U8316 ( .A1(n7807), .A2(n7808), .ZN(n7797) );
  AOI221_X2 U8317 ( .B1(pipeline_regfile_data[114]), .B2(n8247), .C1(
        pipeline_regfile_data[50]), .C2(n8253), .A(n7809), .ZN(n7808) );
  NAND2_X2 U8318 ( .A1(n7810), .A2(n7811), .ZN(n7809) );
  NAND2_X2 U8319 ( .A1(pipeline_regfile_data[242]), .A2(n8255), .ZN(n7811) );
  NAND2_X2 U8320 ( .A1(pipeline_regfile_data[178]), .A2(n8257), .ZN(n7810) );
  AOI221_X2 U8321 ( .B1(pipeline_regfile_data[82]), .B2(n8259), .C1(
        pipeline_regfile_data[18]), .C2(n8262), .A(n7812), .ZN(n7807) );
  NAND2_X2 U8322 ( .A1(n7813), .A2(n7814), .ZN(n7812) );
  NAND2_X2 U8323 ( .A1(pipeline_regfile_data[210]), .A2(n6599), .ZN(n7814) );
  NAND2_X2 U8324 ( .A1(pipeline_regfile_data[146]), .A2(n8271), .ZN(n7813) );
  AOI221_X2 U8325 ( .B1(pipeline_regfile_data[1010]), .B2(n6725), .C1(
        pipeline_regfile_data[754]), .C2(n6721), .A(n7815), .ZN(n7794) );
  INV_X4 U8326 ( .A(n7816), .ZN(n7815) );
  AOI221_X2 U8327 ( .B1(pipeline_regfile_data[562]), .B2(n6726), .C1(
        pipeline_regfile_data[818]), .C2(n6722), .A(n7817), .ZN(n7816) );
  AND2_X1 U8328 ( .A1(pipeline_regfile_data[626]), .A2(n6730), .ZN(n7817) );
  NAND2_X2 U8329 ( .A1(n7819), .A2(n7820), .ZN(n7818) );
  NAND2_X2 U8330 ( .A1(pipeline_regfile_data[658]), .A2(n6731), .ZN(n7820) );
  NAND2_X2 U8331 ( .A1(pipeline_regfile_data[882]), .A2(n6732), .ZN(n7819) );
  AOI221_X2 U8332 ( .B1(pipeline_regfile_data[530]), .B2(n6719), .C1(
        pipeline_regfile_data[978]), .C2(n6723), .A(n7821), .ZN(n7792) );
  INV_X4 U8333 ( .A(n7822), .ZN(n7821) );
  AOI221_X2 U8334 ( .B1(pipeline_regfile_data[786]), .B2(n6727), .C1(
        pipeline_regfile_data[594]), .C2(n6724), .A(n7823), .ZN(n7822) );
  AND2_X1 U8335 ( .A1(pipeline_regfile_data[850]), .A2(n6729), .ZN(n7823) );
  AOI221_X2 U8336 ( .B1(pipeline_regfile_data[947]), .B2(n6728), .C1(
        pipeline_regfile_data[691]), .C2(n6720), .A(n7828), .ZN(n7827) );
  OAI22_X2 U8337 ( .A1(n7829), .A2(n6695), .B1(n7830), .B2(n6663), .ZN(n7828)
         );
  AND2_X1 U8338 ( .A1(n7831), .A2(n7832), .ZN(n7830) );
  AOI221_X2 U8339 ( .B1(pipeline_regfile_data[371]), .B2(n8247), .C1(
        pipeline_regfile_data[307]), .C2(n8253), .A(n7833), .ZN(n7832) );
  NAND2_X2 U8340 ( .A1(n7834), .A2(n7835), .ZN(n7833) );
  NAND2_X2 U8341 ( .A1(pipeline_regfile_data[499]), .A2(n8255), .ZN(n7835) );
  NAND2_X2 U8342 ( .A1(pipeline_regfile_data[435]), .A2(n8257), .ZN(n7834) );
  AOI221_X2 U8343 ( .B1(pipeline_regfile_data[339]), .B2(n8259), .C1(
        pipeline_regfile_data[275]), .C2(n8263), .A(n7836), .ZN(n7831) );
  NAND2_X2 U8344 ( .A1(n7837), .A2(n7838), .ZN(n7836) );
  NAND2_X2 U8345 ( .A1(pipeline_regfile_data[467]), .A2(n6599), .ZN(n7838) );
  NAND2_X2 U8346 ( .A1(pipeline_regfile_data[403]), .A2(n8270), .ZN(n7837) );
  AND2_X1 U8347 ( .A1(n7839), .A2(n7840), .ZN(n7829) );
  AOI221_X2 U8348 ( .B1(pipeline_regfile_data[115]), .B2(n8246), .C1(
        pipeline_regfile_data[51]), .C2(n8252), .A(n7841), .ZN(n7840) );
  NAND2_X2 U8349 ( .A1(n7842), .A2(n7843), .ZN(n7841) );
  NAND2_X2 U8350 ( .A1(pipeline_regfile_data[243]), .A2(n8255), .ZN(n7843) );
  NAND2_X2 U8351 ( .A1(pipeline_regfile_data[179]), .A2(n8257), .ZN(n7842) );
  AOI221_X2 U8352 ( .B1(pipeline_regfile_data[83]), .B2(n8258), .C1(
        pipeline_regfile_data[19]), .C2(n8263), .A(n7844), .ZN(n7839) );
  NAND2_X2 U8353 ( .A1(n7845), .A2(n7846), .ZN(n7844) );
  NAND2_X2 U8354 ( .A1(pipeline_regfile_data[211]), .A2(n6599), .ZN(n7846) );
  NAND2_X2 U8355 ( .A1(pipeline_regfile_data[147]), .A2(n8270), .ZN(n7845) );
  AOI221_X2 U8356 ( .B1(pipeline_regfile_data[1011]), .B2(n6725), .C1(
        pipeline_regfile_data[755]), .C2(n6721), .A(n7847), .ZN(n7826) );
  INV_X4 U8357 ( .A(n7848), .ZN(n7847) );
  AOI221_X2 U8358 ( .B1(pipeline_regfile_data[563]), .B2(n6726), .C1(
        pipeline_regfile_data[819]), .C2(n6722), .A(n7849), .ZN(n7848) );
  AND2_X1 U8359 ( .A1(pipeline_regfile_data[627]), .A2(n6730), .ZN(n7849) );
  NAND2_X2 U8360 ( .A1(n7851), .A2(n7852), .ZN(n7850) );
  NAND2_X2 U8361 ( .A1(pipeline_regfile_data[659]), .A2(n6731), .ZN(n7852) );
  NAND2_X2 U8362 ( .A1(pipeline_regfile_data[883]), .A2(n6732), .ZN(n7851) );
  AOI221_X2 U8363 ( .B1(pipeline_regfile_data[531]), .B2(n6719), .C1(
        pipeline_regfile_data[979]), .C2(n6723), .A(n7853), .ZN(n7824) );
  INV_X4 U8364 ( .A(n7854), .ZN(n7853) );
  AOI221_X2 U8365 ( .B1(pipeline_regfile_data[787]), .B2(n6727), .C1(
        pipeline_regfile_data[595]), .C2(n6724), .A(n7855), .ZN(n7854) );
  AND2_X1 U8366 ( .A1(pipeline_regfile_data[851]), .A2(n6729), .ZN(n7855) );
  AOI221_X2 U8367 ( .B1(pipeline_regfile_data[948]), .B2(n6728), .C1(
        pipeline_regfile_data[692]), .C2(n6720), .A(n7860), .ZN(n7859) );
  OAI22_X2 U8368 ( .A1(n7861), .A2(n6695), .B1(n7862), .B2(n6663), .ZN(n7860)
         );
  AND2_X1 U8369 ( .A1(n7863), .A2(n7864), .ZN(n7862) );
  AOI221_X2 U8370 ( .B1(pipeline_regfile_data[372]), .B2(n8246), .C1(
        pipeline_regfile_data[308]), .C2(n8252), .A(n7865), .ZN(n7864) );
  NAND2_X2 U8371 ( .A1(n7866), .A2(n7867), .ZN(n7865) );
  NAND2_X2 U8372 ( .A1(pipeline_regfile_data[500]), .A2(n8256), .ZN(n7867) );
  NAND2_X2 U8373 ( .A1(pipeline_regfile_data[436]), .A2(n8257), .ZN(n7866) );
  AOI221_X2 U8374 ( .B1(pipeline_regfile_data[340]), .B2(n8258), .C1(
        pipeline_regfile_data[276]), .C2(n8262), .A(n7868), .ZN(n7863) );
  NAND2_X2 U8375 ( .A1(n7869), .A2(n7870), .ZN(n7868) );
  NAND2_X2 U8376 ( .A1(pipeline_regfile_data[468]), .A2(n8268), .ZN(n7870) );
  NAND2_X2 U8377 ( .A1(pipeline_regfile_data[404]), .A2(n8271), .ZN(n7869) );
  AND2_X1 U8378 ( .A1(n7871), .A2(n7872), .ZN(n7861) );
  AOI221_X2 U8379 ( .B1(pipeline_regfile_data[116]), .B2(n8246), .C1(
        pipeline_regfile_data[52]), .C2(n8252), .A(n7873), .ZN(n7872) );
  NAND2_X2 U8380 ( .A1(n7874), .A2(n7875), .ZN(n7873) );
  NAND2_X2 U8381 ( .A1(pipeline_regfile_data[244]), .A2(n8256), .ZN(n7875) );
  NAND2_X2 U8382 ( .A1(pipeline_regfile_data[180]), .A2(n8257), .ZN(n7874) );
  AOI221_X2 U8383 ( .B1(pipeline_regfile_data[84]), .B2(n8258), .C1(
        pipeline_regfile_data[20]), .C2(n8265), .A(n7876), .ZN(n7871) );
  NAND2_X2 U8384 ( .A1(n7877), .A2(n7878), .ZN(n7876) );
  NAND2_X2 U8385 ( .A1(pipeline_regfile_data[212]), .A2(n8268), .ZN(n7878) );
  NAND2_X2 U8386 ( .A1(pipeline_regfile_data[148]), .A2(n8271), .ZN(n7877) );
  AOI221_X2 U8387 ( .B1(pipeline_regfile_data[1012]), .B2(n6725), .C1(
        pipeline_regfile_data[756]), .C2(n6721), .A(n7879), .ZN(n7858) );
  INV_X4 U8388 ( .A(n7880), .ZN(n7879) );
  AOI221_X2 U8389 ( .B1(pipeline_regfile_data[564]), .B2(n6726), .C1(
        pipeline_regfile_data[820]), .C2(n6722), .A(n7881), .ZN(n7880) );
  AND2_X1 U8390 ( .A1(pipeline_regfile_data[628]), .A2(n6730), .ZN(n7881) );
  AOI221_X2 U8391 ( .B1(pipeline_regfile_data[724]), .B2(n6734), .C1(
        pipeline_regfile_data[916]), .C2(n6733), .A(n7882), .ZN(n7857) );
  NAND2_X2 U8392 ( .A1(n7883), .A2(n7884), .ZN(n7882) );
  NAND2_X2 U8393 ( .A1(pipeline_regfile_data[660]), .A2(n6731), .ZN(n7884) );
  NAND2_X2 U8394 ( .A1(pipeline_regfile_data[884]), .A2(n6732), .ZN(n7883) );
  AOI221_X2 U8395 ( .B1(pipeline_regfile_data[532]), .B2(n6719), .C1(
        pipeline_regfile_data[980]), .C2(n6723), .A(n7885), .ZN(n7856) );
  INV_X4 U8396 ( .A(n7886), .ZN(n7885) );
  AOI221_X2 U8397 ( .B1(pipeline_regfile_data[788]), .B2(n6727), .C1(
        pipeline_regfile_data[596]), .C2(n6724), .A(n7887), .ZN(n7886) );
  AND2_X1 U8398 ( .A1(pipeline_regfile_data[852]), .A2(n6729), .ZN(n7887) );
  AOI221_X2 U8399 ( .B1(pipeline_regfile_data[949]), .B2(n6728), .C1(
        pipeline_regfile_data[693]), .C2(n6720), .A(n7892), .ZN(n7891) );
  OAI22_X2 U8400 ( .A1(n7893), .A2(n6695), .B1(n7894), .B2(n6663), .ZN(n7892)
         );
  AND2_X1 U8401 ( .A1(n7895), .A2(n7896), .ZN(n7894) );
  AOI221_X2 U8402 ( .B1(pipeline_regfile_data[373]), .B2(n8246), .C1(
        pipeline_regfile_data[309]), .C2(n8252), .A(n7897), .ZN(n7896) );
  NAND2_X2 U8403 ( .A1(n7898), .A2(n7899), .ZN(n7897) );
  NAND2_X2 U8404 ( .A1(pipeline_regfile_data[501]), .A2(n8256), .ZN(n7899) );
  NAND2_X2 U8405 ( .A1(pipeline_regfile_data[437]), .A2(n8257), .ZN(n7898) );
  AOI221_X2 U8406 ( .B1(pipeline_regfile_data[341]), .B2(n8258), .C1(
        pipeline_regfile_data[277]), .C2(n8265), .A(n7900), .ZN(n7895) );
  NAND2_X2 U8407 ( .A1(n7901), .A2(n7902), .ZN(n7900) );
  NAND2_X2 U8408 ( .A1(pipeline_regfile_data[469]), .A2(n8268), .ZN(n7902) );
  NAND2_X2 U8409 ( .A1(pipeline_regfile_data[405]), .A2(n8270), .ZN(n7901) );
  AND2_X1 U8410 ( .A1(n7903), .A2(n7904), .ZN(n7893) );
  NAND2_X2 U8411 ( .A1(n7906), .A2(n7907), .ZN(n7905) );
  NAND2_X2 U8412 ( .A1(pipeline_regfile_data[245]), .A2(n8256), .ZN(n7907) );
  NAND2_X2 U8413 ( .A1(pipeline_regfile_data[181]), .A2(n8257), .ZN(n7906) );
  AOI221_X2 U8414 ( .B1(pipeline_regfile_data[85]), .B2(n8258), .C1(
        pipeline_regfile_data[21]), .C2(n8262), .A(n7908), .ZN(n7903) );
  NAND2_X2 U8415 ( .A1(n7909), .A2(n7910), .ZN(n7908) );
  NAND2_X2 U8416 ( .A1(pipeline_regfile_data[213]), .A2(n8268), .ZN(n7910) );
  NAND2_X2 U8417 ( .A1(pipeline_regfile_data[149]), .A2(n8271), .ZN(n7909) );
  AOI221_X2 U8418 ( .B1(pipeline_regfile_data[1013]), .B2(n6725), .C1(
        pipeline_regfile_data[757]), .C2(n6721), .A(n7911), .ZN(n7890) );
  INV_X4 U8419 ( .A(n7912), .ZN(n7911) );
  AOI221_X2 U8420 ( .B1(pipeline_regfile_data[565]), .B2(n6726), .C1(
        pipeline_regfile_data[821]), .C2(n6722), .A(n7913), .ZN(n7912) );
  AND2_X1 U8421 ( .A1(pipeline_regfile_data[629]), .A2(n6730), .ZN(n7913) );
  NAND2_X2 U8422 ( .A1(n7915), .A2(n7916), .ZN(n7914) );
  NAND2_X2 U8423 ( .A1(pipeline_regfile_data[661]), .A2(n6731), .ZN(n7916) );
  NAND2_X2 U8424 ( .A1(pipeline_regfile_data[885]), .A2(n6732), .ZN(n7915) );
  AOI221_X2 U8425 ( .B1(pipeline_regfile_data[533]), .B2(n6719), .C1(
        pipeline_regfile_data[981]), .C2(n6723), .A(n7917), .ZN(n7888) );
  INV_X4 U8426 ( .A(n7918), .ZN(n7917) );
  AOI221_X2 U8427 ( .B1(pipeline_regfile_data[789]), .B2(n6727), .C1(
        pipeline_regfile_data[597]), .C2(n6724), .A(n7919), .ZN(n7918) );
  AND2_X1 U8428 ( .A1(pipeline_regfile_data[853]), .A2(n6729), .ZN(n7919) );
  AOI221_X2 U8429 ( .B1(pipeline_regfile_data[950]), .B2(n6728), .C1(
        pipeline_regfile_data[694]), .C2(n6720), .A(n7924), .ZN(n7923) );
  OAI22_X2 U8430 ( .A1(n7925), .A2(n6695), .B1(n7926), .B2(n6663), .ZN(n7924)
         );
  AND2_X1 U8431 ( .A1(n7927), .A2(n7928), .ZN(n7926) );
  AOI221_X2 U8432 ( .B1(pipeline_regfile_data[374]), .B2(n8246), .C1(
        pipeline_regfile_data[310]), .C2(n8252), .A(n7929), .ZN(n7928) );
  NAND2_X2 U8433 ( .A1(n7930), .A2(n7931), .ZN(n7929) );
  NAND2_X2 U8434 ( .A1(pipeline_regfile_data[502]), .A2(n8256), .ZN(n7931) );
  NAND2_X2 U8435 ( .A1(pipeline_regfile_data[438]), .A2(n8257), .ZN(n7930) );
  AOI221_X2 U8436 ( .B1(pipeline_regfile_data[342]), .B2(n8258), .C1(
        pipeline_regfile_data[278]), .C2(n8262), .A(n7932), .ZN(n7927) );
  NAND2_X2 U8437 ( .A1(n7933), .A2(n7934), .ZN(n7932) );
  NAND2_X2 U8438 ( .A1(pipeline_regfile_data[470]), .A2(n8268), .ZN(n7934) );
  NAND2_X2 U8439 ( .A1(pipeline_regfile_data[406]), .A2(n8269), .ZN(n7933) );
  AND2_X1 U8440 ( .A1(n7935), .A2(n7936), .ZN(n7925) );
  NAND2_X2 U8441 ( .A1(n7938), .A2(n7939), .ZN(n7937) );
  NAND2_X2 U8442 ( .A1(pipeline_regfile_data[246]), .A2(n8256), .ZN(n7939) );
  NAND2_X2 U8443 ( .A1(pipeline_regfile_data[182]), .A2(n8257), .ZN(n7938) );
  AOI221_X2 U8444 ( .B1(pipeline_regfile_data[86]), .B2(n8258), .C1(
        pipeline_regfile_data[22]), .C2(n8265), .A(n7940), .ZN(n7935) );
  NAND2_X2 U8445 ( .A1(n7941), .A2(n7942), .ZN(n7940) );
  NAND2_X2 U8446 ( .A1(pipeline_regfile_data[214]), .A2(n8268), .ZN(n7942) );
  NAND2_X2 U8447 ( .A1(pipeline_regfile_data[150]), .A2(n8271), .ZN(n7941) );
  AOI221_X2 U8448 ( .B1(pipeline_regfile_data[1014]), .B2(n6725), .C1(
        pipeline_regfile_data[758]), .C2(n6721), .A(n7943), .ZN(n7922) );
  INV_X4 U8449 ( .A(n7944), .ZN(n7943) );
  AOI221_X2 U8450 ( .B1(pipeline_regfile_data[566]), .B2(n6726), .C1(
        pipeline_regfile_data[822]), .C2(n6722), .A(n7945), .ZN(n7944) );
  AND2_X1 U8451 ( .A1(pipeline_regfile_data[630]), .A2(n6730), .ZN(n7945) );
  NAND2_X2 U8452 ( .A1(n7947), .A2(n7948), .ZN(n7946) );
  NAND2_X2 U8453 ( .A1(pipeline_regfile_data[662]), .A2(n6731), .ZN(n7948) );
  NAND2_X2 U8454 ( .A1(pipeline_regfile_data[886]), .A2(n6732), .ZN(n7947) );
  AOI221_X2 U8455 ( .B1(pipeline_regfile_data[534]), .B2(n6719), .C1(
        pipeline_regfile_data[982]), .C2(n6723), .A(n7949), .ZN(n7920) );
  INV_X4 U8456 ( .A(n7950), .ZN(n7949) );
  AOI221_X2 U8457 ( .B1(pipeline_regfile_data[790]), .B2(n6727), .C1(
        pipeline_regfile_data[598]), .C2(n6724), .A(n7951), .ZN(n7950) );
  AND2_X1 U8458 ( .A1(pipeline_regfile_data[854]), .A2(n6729), .ZN(n7951) );
  AOI221_X2 U8459 ( .B1(pipeline_regfile_data[951]), .B2(n6728), .C1(
        pipeline_regfile_data[695]), .C2(n6720), .A(n7956), .ZN(n7955) );
  OAI22_X2 U8460 ( .A1(n7957), .A2(n6695), .B1(n7958), .B2(n6663), .ZN(n7956)
         );
  AND2_X1 U8461 ( .A1(n7959), .A2(n7960), .ZN(n7958) );
  AOI221_X2 U8462 ( .B1(pipeline_regfile_data[375]), .B2(n8246), .C1(
        pipeline_regfile_data[311]), .C2(n8252), .A(n7961), .ZN(n7960) );
  NAND2_X2 U8463 ( .A1(n7962), .A2(n7963), .ZN(n7961) );
  NAND2_X2 U8464 ( .A1(pipeline_regfile_data[503]), .A2(n8256), .ZN(n7963) );
  NAND2_X2 U8465 ( .A1(pipeline_regfile_data[439]), .A2(n8257), .ZN(n7962) );
  AOI221_X2 U8466 ( .B1(pipeline_regfile_data[343]), .B2(n8258), .C1(
        pipeline_regfile_data[279]), .C2(n8265), .A(n7964), .ZN(n7959) );
  NAND2_X2 U8467 ( .A1(n7965), .A2(n7966), .ZN(n7964) );
  NAND2_X2 U8468 ( .A1(pipeline_regfile_data[471]), .A2(n8268), .ZN(n7966) );
  NAND2_X2 U8469 ( .A1(pipeline_regfile_data[407]), .A2(n8270), .ZN(n7965) );
  AND2_X1 U8470 ( .A1(n7967), .A2(n7968), .ZN(n7957) );
  AOI221_X2 U8471 ( .B1(pipeline_regfile_data[119]), .B2(n8246), .C1(
        pipeline_regfile_data[55]), .C2(n8252), .A(n7969), .ZN(n7968) );
  NAND2_X2 U8472 ( .A1(n7970), .A2(n7971), .ZN(n7969) );
  NAND2_X2 U8473 ( .A1(pipeline_regfile_data[247]), .A2(n8256), .ZN(n7971) );
  NAND2_X2 U8474 ( .A1(pipeline_regfile_data[183]), .A2(n8257), .ZN(n7970) );
  AOI221_X2 U8475 ( .B1(pipeline_regfile_data[87]), .B2(n8258), .C1(
        pipeline_regfile_data[23]), .C2(n8265), .A(n7972), .ZN(n7967) );
  NAND2_X2 U8476 ( .A1(n7973), .A2(n7974), .ZN(n7972) );
  NAND2_X2 U8477 ( .A1(pipeline_regfile_data[215]), .A2(n8268), .ZN(n7974) );
  NAND2_X2 U8478 ( .A1(pipeline_regfile_data[151]), .A2(n8269), .ZN(n7973) );
  AOI221_X2 U8479 ( .B1(pipeline_regfile_data[1015]), .B2(n6725), .C1(
        pipeline_regfile_data[759]), .C2(n6721), .A(n7975), .ZN(n7954) );
  INV_X4 U8480 ( .A(n7976), .ZN(n7975) );
  AOI221_X2 U8481 ( .B1(pipeline_regfile_data[567]), .B2(n6726), .C1(
        pipeline_regfile_data[823]), .C2(n6722), .A(n7977), .ZN(n7976) );
  AND2_X1 U8482 ( .A1(pipeline_regfile_data[631]), .A2(n6730), .ZN(n7977) );
  NAND2_X2 U8483 ( .A1(n7979), .A2(n7980), .ZN(n7978) );
  NAND2_X2 U8484 ( .A1(pipeline_regfile_data[663]), .A2(n6731), .ZN(n7980) );
  NAND2_X2 U8485 ( .A1(pipeline_regfile_data[887]), .A2(n6732), .ZN(n7979) );
  AOI221_X2 U8486 ( .B1(pipeline_regfile_data[535]), .B2(n6719), .C1(
        pipeline_regfile_data[983]), .C2(n6723), .A(n7981), .ZN(n7952) );
  INV_X4 U8487 ( .A(n7982), .ZN(n7981) );
  AOI221_X2 U8488 ( .B1(pipeline_regfile_data[791]), .B2(n6727), .C1(
        pipeline_regfile_data[599]), .C2(n6724), .A(n7983), .ZN(n7982) );
  AND2_X1 U8489 ( .A1(pipeline_regfile_data[855]), .A2(n6729), .ZN(n7983) );
  OAI22_X2 U8490 ( .A1(n7989), .A2(n6695), .B1(n7990), .B2(n6663), .ZN(n7988)
         );
  AND2_X1 U8491 ( .A1(n7991), .A2(n7992), .ZN(n7990) );
  AOI221_X2 U8492 ( .B1(pipeline_regfile_data[376]), .B2(n8246), .C1(
        pipeline_regfile_data[312]), .C2(n8252), .A(n7993), .ZN(n7992) );
  NAND2_X2 U8493 ( .A1(n7994), .A2(n7995), .ZN(n7993) );
  NAND2_X2 U8494 ( .A1(pipeline_regfile_data[504]), .A2(n8256), .ZN(n7995) );
  NAND2_X2 U8495 ( .A1(pipeline_regfile_data[440]), .A2(n8257), .ZN(n7994) );
  AOI221_X2 U8496 ( .B1(pipeline_regfile_data[344]), .B2(n8258), .C1(
        pipeline_regfile_data[280]), .C2(n8264), .A(n7996), .ZN(n7991) );
  NAND2_X2 U8497 ( .A1(n7997), .A2(n7998), .ZN(n7996) );
  NAND2_X2 U8498 ( .A1(pipeline_regfile_data[472]), .A2(n8268), .ZN(n7998) );
  NAND2_X2 U8499 ( .A1(pipeline_regfile_data[408]), .A2(n8271), .ZN(n7997) );
  AND2_X1 U8500 ( .A1(n7999), .A2(n8000), .ZN(n7989) );
  AOI221_X2 U8501 ( .B1(pipeline_regfile_data[120]), .B2(n8246), .C1(
        pipeline_regfile_data[56]), .C2(n8252), .A(n8001), .ZN(n8000) );
  NAND2_X2 U8502 ( .A1(n8002), .A2(n8003), .ZN(n8001) );
  NAND2_X2 U8503 ( .A1(pipeline_regfile_data[248]), .A2(n8256), .ZN(n8003) );
  NAND2_X2 U8504 ( .A1(pipeline_regfile_data[184]), .A2(n8257), .ZN(n8002) );
  AOI221_X2 U8505 ( .B1(pipeline_regfile_data[88]), .B2(n8258), .C1(
        pipeline_regfile_data[24]), .C2(n8265), .A(n8004), .ZN(n7999) );
  NAND2_X2 U8506 ( .A1(n8005), .A2(n8006), .ZN(n8004) );
  NAND2_X2 U8507 ( .A1(pipeline_regfile_data[216]), .A2(n8268), .ZN(n8006) );
  NAND2_X2 U8508 ( .A1(pipeline_regfile_data[152]), .A2(n8271), .ZN(n8005) );
  AOI221_X2 U8509 ( .B1(pipeline_regfile_data[1016]), .B2(n6725), .C1(
        pipeline_regfile_data[760]), .C2(n6721), .A(n8007), .ZN(n7986) );
  INV_X4 U8510 ( .A(n8008), .ZN(n8007) );
  AOI221_X2 U8511 ( .B1(pipeline_regfile_data[568]), .B2(n6726), .C1(
        pipeline_regfile_data[824]), .C2(n6722), .A(n8009), .ZN(n8008) );
  AND2_X1 U8512 ( .A1(pipeline_regfile_data[632]), .A2(n6730), .ZN(n8009) );
  AOI221_X2 U8513 ( .B1(pipeline_regfile_data[728]), .B2(n6734), .C1(
        pipeline_regfile_data[920]), .C2(n6733), .A(n8010), .ZN(n7985) );
  NAND2_X2 U8514 ( .A1(n8011), .A2(n8012), .ZN(n8010) );
  NAND2_X2 U8515 ( .A1(pipeline_regfile_data[664]), .A2(n6731), .ZN(n8012) );
  NAND2_X2 U8516 ( .A1(pipeline_regfile_data[888]), .A2(n6732), .ZN(n8011) );
  AOI221_X2 U8517 ( .B1(pipeline_regfile_data[536]), .B2(n6719), .C1(
        pipeline_regfile_data[984]), .C2(n6723), .A(n8013), .ZN(n7984) );
  INV_X4 U8518 ( .A(n8014), .ZN(n8013) );
  AOI221_X2 U8519 ( .B1(pipeline_regfile_data[792]), .B2(n6727), .C1(
        pipeline_regfile_data[600]), .C2(n6724), .A(n8015), .ZN(n8014) );
  AND2_X1 U8520 ( .A1(pipeline_regfile_data[856]), .A2(n6729), .ZN(n8015) );
  AOI221_X2 U8521 ( .B1(pipeline_regfile_data[953]), .B2(n6728), .C1(
        pipeline_regfile_data[697]), .C2(n6720), .A(n8020), .ZN(n8019) );
  OAI22_X2 U8522 ( .A1(n8021), .A2(n6695), .B1(n8022), .B2(n6663), .ZN(n8020)
         );
  AND2_X1 U8523 ( .A1(n8023), .A2(n8024), .ZN(n8022) );
  AOI221_X2 U8524 ( .B1(pipeline_regfile_data[377]), .B2(n8246), .C1(
        pipeline_regfile_data[313]), .C2(n8252), .A(n8025), .ZN(n8024) );
  NAND2_X2 U8525 ( .A1(n8026), .A2(n8027), .ZN(n8025) );
  NAND2_X2 U8526 ( .A1(pipeline_regfile_data[505]), .A2(n8256), .ZN(n8027) );
  NAND2_X2 U8527 ( .A1(pipeline_regfile_data[441]), .A2(n8257), .ZN(n8026) );
  AOI221_X2 U8528 ( .B1(pipeline_regfile_data[345]), .B2(n8258), .C1(
        pipeline_regfile_data[281]), .C2(n8263), .A(n8028), .ZN(n8023) );
  NAND2_X2 U8529 ( .A1(n8029), .A2(n8030), .ZN(n8028) );
  NAND2_X2 U8530 ( .A1(pipeline_regfile_data[473]), .A2(n8268), .ZN(n8030) );
  NAND2_X2 U8531 ( .A1(pipeline_regfile_data[409]), .A2(n8270), .ZN(n8029) );
  AND2_X1 U8532 ( .A1(n8031), .A2(n8032), .ZN(n8021) );
  NAND2_X2 U8533 ( .A1(n8034), .A2(n8035), .ZN(n8033) );
  NAND2_X2 U8534 ( .A1(pipeline_regfile_data[249]), .A2(n8256), .ZN(n8035) );
  NAND2_X2 U8535 ( .A1(pipeline_regfile_data[185]), .A2(n8257), .ZN(n8034) );
  AOI221_X2 U8536 ( .B1(pipeline_regfile_data[89]), .B2(n8258), .C1(
        pipeline_regfile_data[25]), .C2(n8262), .A(n8036), .ZN(n8031) );
  NAND2_X2 U8537 ( .A1(n8037), .A2(n8038), .ZN(n8036) );
  NAND2_X2 U8538 ( .A1(pipeline_regfile_data[217]), .A2(n8268), .ZN(n8038) );
  NAND2_X2 U8539 ( .A1(pipeline_regfile_data[153]), .A2(n8270), .ZN(n8037) );
  AOI221_X2 U8540 ( .B1(pipeline_regfile_data[1017]), .B2(n6725), .C1(
        pipeline_regfile_data[761]), .C2(n6721), .A(n8039), .ZN(n8018) );
  INV_X4 U8541 ( .A(n8040), .ZN(n8039) );
  AOI221_X2 U8542 ( .B1(pipeline_regfile_data[569]), .B2(n6726), .C1(
        pipeline_regfile_data[825]), .C2(n6722), .A(n8041), .ZN(n8040) );
  AND2_X1 U8543 ( .A1(pipeline_regfile_data[633]), .A2(n6730), .ZN(n8041) );
  NAND2_X2 U8544 ( .A1(n8043), .A2(n8044), .ZN(n8042) );
  NAND2_X2 U8545 ( .A1(pipeline_regfile_data[665]), .A2(n6731), .ZN(n8044) );
  NAND2_X2 U8546 ( .A1(pipeline_regfile_data[889]), .A2(n6732), .ZN(n8043) );
  AOI221_X2 U8547 ( .B1(pipeline_regfile_data[537]), .B2(n6719), .C1(
        pipeline_regfile_data[985]), .C2(n6723), .A(n8045), .ZN(n8016) );
  INV_X4 U8548 ( .A(n8046), .ZN(n8045) );
  AOI221_X2 U8549 ( .B1(pipeline_regfile_data[793]), .B2(n6727), .C1(
        pipeline_regfile_data[601]), .C2(n6724), .A(n8047), .ZN(n8046) );
  AND2_X1 U8550 ( .A1(pipeline_regfile_data[857]), .A2(n6729), .ZN(n8047) );
  OAI22_X2 U8551 ( .A1(n8052), .A2(n6695), .B1(n8053), .B2(n6663), .ZN(n8051)
         );
  AND2_X1 U8552 ( .A1(n8054), .A2(n8055), .ZN(n8053) );
  AOI221_X2 U8553 ( .B1(pipeline_regfile_data[378]), .B2(n8249), .C1(
        pipeline_regfile_data[314]), .C2(n8251), .A(n8056), .ZN(n8055) );
  NAND2_X2 U8554 ( .A1(n8057), .A2(n8058), .ZN(n8056) );
  NAND2_X2 U8555 ( .A1(pipeline_regfile_data[506]), .A2(n8256), .ZN(n8058) );
  NAND2_X2 U8556 ( .A1(pipeline_regfile_data[442]), .A2(n8257), .ZN(n8057) );
  AOI221_X2 U8557 ( .B1(pipeline_regfile_data[346]), .B2(n8261), .C1(
        pipeline_regfile_data[282]), .C2(n8265), .A(n8059), .ZN(n8054) );
  NAND2_X2 U8558 ( .A1(n8060), .A2(n8061), .ZN(n8059) );
  NAND2_X2 U8559 ( .A1(pipeline_regfile_data[474]), .A2(n8268), .ZN(n8061) );
  NAND2_X2 U8560 ( .A1(pipeline_regfile_data[410]), .A2(n8271), .ZN(n8060) );
  AND2_X1 U8561 ( .A1(n8062), .A2(n8063), .ZN(n8052) );
  AOI221_X2 U8562 ( .B1(pipeline_regfile_data[122]), .B2(n8247), .C1(
        pipeline_regfile_data[58]), .C2(n8251), .A(n8064), .ZN(n8063) );
  NAND2_X2 U8563 ( .A1(n8065), .A2(n8066), .ZN(n8064) );
  NAND2_X2 U8564 ( .A1(pipeline_regfile_data[250]), .A2(n8256), .ZN(n8066) );
  NAND2_X2 U8565 ( .A1(pipeline_regfile_data[186]), .A2(n8257), .ZN(n8065) );
  AOI221_X2 U8566 ( .B1(pipeline_regfile_data[90]), .B2(n8261), .C1(
        pipeline_regfile_data[26]), .C2(n8263), .A(n8067), .ZN(n8062) );
  NAND2_X2 U8567 ( .A1(n8068), .A2(n8069), .ZN(n8067) );
  NAND2_X2 U8568 ( .A1(pipeline_regfile_data[218]), .A2(n8268), .ZN(n8069) );
  NAND2_X2 U8569 ( .A1(pipeline_regfile_data[154]), .A2(n8269), .ZN(n8068) );
  AOI221_X2 U8570 ( .B1(pipeline_regfile_data[1018]), .B2(n6725), .C1(
        pipeline_regfile_data[762]), .C2(n6721), .A(n8070), .ZN(n8050) );
  INV_X4 U8571 ( .A(n8071), .ZN(n8070) );
  AOI221_X2 U8572 ( .B1(pipeline_regfile_data[570]), .B2(n6726), .C1(
        pipeline_regfile_data[826]), .C2(n6722), .A(n8072), .ZN(n8071) );
  AND2_X1 U8573 ( .A1(pipeline_regfile_data[634]), .A2(n6730), .ZN(n8072) );
  AOI221_X2 U8574 ( .B1(pipeline_regfile_data[730]), .B2(n6734), .C1(
        pipeline_regfile_data[922]), .C2(n6733), .A(n8073), .ZN(n8049) );
  NAND2_X2 U8575 ( .A1(n8074), .A2(n8075), .ZN(n8073) );
  NAND2_X2 U8576 ( .A1(pipeline_regfile_data[666]), .A2(n6731), .ZN(n8075) );
  NAND2_X2 U8577 ( .A1(pipeline_regfile_data[890]), .A2(n6732), .ZN(n8074) );
  AOI221_X2 U8578 ( .B1(pipeline_regfile_data[538]), .B2(n6719), .C1(
        pipeline_regfile_data[986]), .C2(n6723), .A(n8076), .ZN(n8048) );
  INV_X4 U8579 ( .A(n8077), .ZN(n8076) );
  AOI221_X2 U8580 ( .B1(pipeline_regfile_data[794]), .B2(n6727), .C1(
        pipeline_regfile_data[602]), .C2(n6724), .A(n8078), .ZN(n8077) );
  AND2_X1 U8581 ( .A1(pipeline_regfile_data[858]), .A2(n6729), .ZN(n8078) );
  OAI22_X2 U8582 ( .A1(n8084), .A2(n6695), .B1(n8085), .B2(n6663), .ZN(n8083)
         );
  AOI221_X2 U8583 ( .B1(pipeline_regfile_data[379]), .B2(n8246), .C1(
        pipeline_regfile_data[315]), .C2(n8251), .A(n8088), .ZN(n8087) );
  NAND2_X2 U8584 ( .A1(n8089), .A2(n8090), .ZN(n8088) );
  NAND2_X2 U8585 ( .A1(pipeline_regfile_data[507]), .A2(n8256), .ZN(n8090) );
  NAND2_X2 U8586 ( .A1(pipeline_regfile_data[443]), .A2(n8257), .ZN(n8089) );
  AOI221_X2 U8587 ( .B1(pipeline_regfile_data[347]), .B2(n8259), .C1(
        pipeline_regfile_data[283]), .C2(n8263), .A(n8091), .ZN(n8086) );
  NAND2_X2 U8588 ( .A1(n8092), .A2(n8093), .ZN(n8091) );
  NAND2_X2 U8589 ( .A1(pipeline_regfile_data[475]), .A2(n8268), .ZN(n8093) );
  NAND2_X2 U8590 ( .A1(pipeline_regfile_data[411]), .A2(n8270), .ZN(n8092) );
  AND2_X1 U8591 ( .A1(n8094), .A2(n8095), .ZN(n8084) );
  AOI221_X2 U8592 ( .B1(pipeline_regfile_data[123]), .B2(n8249), .C1(
        pipeline_regfile_data[59]), .C2(n8251), .A(n8096), .ZN(n8095) );
  NAND2_X2 U8593 ( .A1(n8097), .A2(n8098), .ZN(n8096) );
  NAND2_X2 U8594 ( .A1(pipeline_regfile_data[251]), .A2(n8255), .ZN(n8098) );
  NAND2_X2 U8595 ( .A1(pipeline_regfile_data[187]), .A2(n8257), .ZN(n8097) );
  AOI221_X2 U8596 ( .B1(pipeline_regfile_data[91]), .B2(n8261), .C1(
        pipeline_regfile_data[27]), .C2(n8265), .A(n8099), .ZN(n8094) );
  NAND2_X2 U8597 ( .A1(n8100), .A2(n8101), .ZN(n8099) );
  NAND2_X2 U8598 ( .A1(pipeline_regfile_data[219]), .A2(n6599), .ZN(n8101) );
  NAND2_X2 U8599 ( .A1(pipeline_regfile_data[155]), .A2(n8270), .ZN(n8100) );
  AOI221_X2 U8600 ( .B1(pipeline_regfile_data[1019]), .B2(n6725), .C1(
        pipeline_regfile_data[763]), .C2(n6721), .A(n8102), .ZN(n8081) );
  INV_X4 U8601 ( .A(n8103), .ZN(n8102) );
  AOI221_X2 U8602 ( .B1(pipeline_regfile_data[571]), .B2(n6726), .C1(
        pipeline_regfile_data[827]), .C2(n6722), .A(n8104), .ZN(n8103) );
  AND2_X1 U8603 ( .A1(pipeline_regfile_data[635]), .A2(n6730), .ZN(n8104) );
  NAND2_X2 U8604 ( .A1(n8106), .A2(n8107), .ZN(n8105) );
  NAND2_X2 U8605 ( .A1(pipeline_regfile_data[667]), .A2(n6731), .ZN(n8107) );
  NAND2_X2 U8606 ( .A1(pipeline_regfile_data[891]), .A2(n6732), .ZN(n8106) );
  AOI221_X2 U8607 ( .B1(pipeline_regfile_data[539]), .B2(n6719), .C1(
        pipeline_regfile_data[987]), .C2(n6723), .A(n8108), .ZN(n8079) );
  INV_X4 U8608 ( .A(n8109), .ZN(n8108) );
  AOI221_X2 U8609 ( .B1(pipeline_regfile_data[795]), .B2(n6727), .C1(
        pipeline_regfile_data[603]), .C2(n6724), .A(n8110), .ZN(n8109) );
  AND2_X1 U8610 ( .A1(pipeline_regfile_data[859]), .A2(n6729), .ZN(n8110) );
  AOI221_X2 U8611 ( .B1(pipeline_regfile_data[956]), .B2(n6728), .C1(
        pipeline_regfile_data[700]), .C2(n6720), .A(n8115), .ZN(n8114) );
  OAI22_X2 U8612 ( .A1(n8116), .A2(n6695), .B1(n8117), .B2(n6663), .ZN(n8115)
         );
  AND2_X1 U8613 ( .A1(n8118), .A2(n8119), .ZN(n8117) );
  AOI221_X2 U8614 ( .B1(pipeline_regfile_data[380]), .B2(n8249), .C1(
        pipeline_regfile_data[316]), .C2(n8251), .A(n8120), .ZN(n8119) );
  NAND2_X2 U8615 ( .A1(n8121), .A2(n8122), .ZN(n8120) );
  NAND2_X2 U8616 ( .A1(pipeline_regfile_data[508]), .A2(n8256), .ZN(n8122) );
  NAND2_X2 U8617 ( .A1(pipeline_regfile_data[444]), .A2(n8257), .ZN(n8121) );
  AOI221_X2 U8618 ( .B1(pipeline_regfile_data[348]), .B2(n8261), .C1(
        pipeline_regfile_data[284]), .C2(n8263), .A(n8123), .ZN(n8118) );
  NAND2_X2 U8619 ( .A1(n8124), .A2(n8125), .ZN(n8123) );
  NAND2_X2 U8620 ( .A1(pipeline_regfile_data[476]), .A2(n8268), .ZN(n8125) );
  NAND2_X2 U8621 ( .A1(pipeline_regfile_data[412]), .A2(n8270), .ZN(n8124) );
  AND2_X1 U8622 ( .A1(n8126), .A2(n8127), .ZN(n8116) );
  AOI221_X2 U8623 ( .B1(pipeline_regfile_data[124]), .B2(n8249), .C1(
        pipeline_regfile_data[60]), .C2(n8251), .A(n8128), .ZN(n8127) );
  NAND2_X2 U8624 ( .A1(n8129), .A2(n8130), .ZN(n8128) );
  NAND2_X2 U8625 ( .A1(pipeline_regfile_data[252]), .A2(n8255), .ZN(n8130) );
  NAND2_X2 U8626 ( .A1(pipeline_regfile_data[188]), .A2(n8257), .ZN(n8129) );
  AOI221_X2 U8627 ( .B1(pipeline_regfile_data[92]), .B2(n8261), .C1(
        pipeline_regfile_data[28]), .C2(n8264), .A(n8131), .ZN(n8126) );
  NAND2_X2 U8628 ( .A1(n8132), .A2(n8133), .ZN(n8131) );
  NAND2_X2 U8629 ( .A1(pipeline_regfile_data[220]), .A2(n6599), .ZN(n8133) );
  NAND2_X2 U8630 ( .A1(pipeline_regfile_data[156]), .A2(n8271), .ZN(n8132) );
  AOI221_X2 U8631 ( .B1(pipeline_regfile_data[1020]), .B2(n6725), .C1(
        pipeline_regfile_data[764]), .C2(n6721), .A(n8134), .ZN(n8113) );
  INV_X4 U8632 ( .A(n8135), .ZN(n8134) );
  AOI221_X2 U8633 ( .B1(pipeline_regfile_data[572]), .B2(n6726), .C1(
        pipeline_regfile_data[828]), .C2(n6722), .A(n8136), .ZN(n8135) );
  AND2_X1 U8634 ( .A1(pipeline_regfile_data[636]), .A2(n6730), .ZN(n8136) );
  NAND2_X2 U8635 ( .A1(n8138), .A2(n8139), .ZN(n8137) );
  NAND2_X2 U8636 ( .A1(pipeline_regfile_data[668]), .A2(n6731), .ZN(n8139) );
  NAND2_X2 U8637 ( .A1(pipeline_regfile_data[892]), .A2(n6732), .ZN(n8138) );
  AOI221_X2 U8638 ( .B1(pipeline_regfile_data[540]), .B2(n6719), .C1(
        pipeline_regfile_data[988]), .C2(n6723), .A(n8140), .ZN(n8111) );
  INV_X4 U8639 ( .A(n8141), .ZN(n8140) );
  AOI221_X2 U8640 ( .B1(pipeline_regfile_data[796]), .B2(n6727), .C1(
        pipeline_regfile_data[604]), .C2(n6724), .A(n8142), .ZN(n8141) );
  AND2_X1 U8641 ( .A1(pipeline_regfile_data[860]), .A2(n6729), .ZN(n8142) );
  AOI221_X2 U8642 ( .B1(pipeline_regfile_data[957]), .B2(n6728), .C1(
        pipeline_regfile_data[701]), .C2(n6720), .A(n8147), .ZN(n8146) );
  OAI22_X2 U8643 ( .A1(n8148), .A2(n6695), .B1(n8149), .B2(n6663), .ZN(n8147)
         );
  AND2_X1 U8644 ( .A1(n8150), .A2(n8151), .ZN(n8149) );
  AOI221_X2 U8645 ( .B1(pipeline_regfile_data[381]), .B2(n8247), .C1(
        pipeline_regfile_data[317]), .C2(n8251), .A(n8152), .ZN(n8151) );
  NAND2_X2 U8646 ( .A1(n8153), .A2(n8154), .ZN(n8152) );
  NAND2_X2 U8647 ( .A1(pipeline_regfile_data[509]), .A2(n8255), .ZN(n8154) );
  NAND2_X2 U8648 ( .A1(pipeline_regfile_data[445]), .A2(n8257), .ZN(n8153) );
  AOI221_X2 U8649 ( .B1(pipeline_regfile_data[349]), .B2(n8259), .C1(
        pipeline_regfile_data[285]), .C2(n8263), .A(n8155), .ZN(n8150) );
  NAND2_X2 U8650 ( .A1(n8156), .A2(n8157), .ZN(n8155) );
  NAND2_X2 U8651 ( .A1(pipeline_regfile_data[477]), .A2(n6599), .ZN(n8157) );
  NAND2_X2 U8652 ( .A1(pipeline_regfile_data[413]), .A2(n8269), .ZN(n8156) );
  AND2_X1 U8653 ( .A1(n8158), .A2(n8159), .ZN(n8148) );
  AOI221_X2 U8654 ( .B1(pipeline_regfile_data[125]), .B2(n8249), .C1(
        pipeline_regfile_data[61]), .C2(n8251), .A(n8160), .ZN(n8159) );
  NAND2_X2 U8655 ( .A1(n8161), .A2(n8162), .ZN(n8160) );
  NAND2_X2 U8656 ( .A1(pipeline_regfile_data[253]), .A2(n8255), .ZN(n8162) );
  NAND2_X2 U8657 ( .A1(pipeline_regfile_data[189]), .A2(n8257), .ZN(n8161) );
  AOI221_X2 U8658 ( .B1(pipeline_regfile_data[93]), .B2(n8261), .C1(
        pipeline_regfile_data[29]), .C2(n8264), .A(n8163), .ZN(n8158) );
  NAND2_X2 U8659 ( .A1(n8164), .A2(n8165), .ZN(n8163) );
  NAND2_X2 U8660 ( .A1(pipeline_regfile_data[221]), .A2(n6599), .ZN(n8165) );
  NAND2_X2 U8661 ( .A1(pipeline_regfile_data[157]), .A2(n8269), .ZN(n8164) );
  AOI221_X2 U8662 ( .B1(pipeline_regfile_data[1021]), .B2(n6725), .C1(
        pipeline_regfile_data[765]), .C2(n6721), .A(n8166), .ZN(n8145) );
  INV_X4 U8663 ( .A(n8167), .ZN(n8166) );
  AOI221_X2 U8664 ( .B1(pipeline_regfile_data[573]), .B2(n6726), .C1(
        pipeline_regfile_data[829]), .C2(n6722), .A(n8168), .ZN(n8167) );
  AND2_X1 U8665 ( .A1(pipeline_regfile_data[637]), .A2(n6730), .ZN(n8168) );
  NAND2_X2 U8666 ( .A1(n8170), .A2(n8171), .ZN(n8169) );
  NAND2_X2 U8667 ( .A1(pipeline_regfile_data[669]), .A2(n6731), .ZN(n8171) );
  NAND2_X2 U8668 ( .A1(pipeline_regfile_data[893]), .A2(n6732), .ZN(n8170) );
  AOI221_X2 U8669 ( .B1(pipeline_regfile_data[541]), .B2(n6719), .C1(
        pipeline_regfile_data[989]), .C2(n6723), .A(n8172), .ZN(n8143) );
  INV_X4 U8670 ( .A(n8173), .ZN(n8172) );
  AOI221_X2 U8671 ( .B1(pipeline_regfile_data[797]), .B2(n6727), .C1(
        pipeline_regfile_data[605]), .C2(n6724), .A(n8174), .ZN(n8173) );
  AND2_X1 U8672 ( .A1(pipeline_regfile_data[861]), .A2(n6729), .ZN(n8174) );
  AOI221_X2 U8673 ( .B1(pipeline_regfile_data[958]), .B2(n6728), .C1(
        pipeline_regfile_data[702]), .C2(n6720), .A(n8179), .ZN(n8178) );
  OAI22_X2 U8674 ( .A1(n8180), .A2(n6695), .B1(n8181), .B2(n6663), .ZN(n8179)
         );
  AND2_X1 U8675 ( .A1(n8182), .A2(n8183), .ZN(n8181) );
  AOI221_X2 U8676 ( .B1(pipeline_regfile_data[382]), .B2(n8249), .C1(
        pipeline_regfile_data[318]), .C2(n8251), .A(n8184), .ZN(n8183) );
  NAND2_X2 U8677 ( .A1(n8185), .A2(n8186), .ZN(n8184) );
  NAND2_X2 U8678 ( .A1(pipeline_regfile_data[510]), .A2(n8255), .ZN(n8186) );
  NAND2_X2 U8679 ( .A1(pipeline_regfile_data[446]), .A2(n8257), .ZN(n8185) );
  AOI221_X2 U8680 ( .B1(pipeline_regfile_data[350]), .B2(n8261), .C1(
        pipeline_regfile_data[286]), .C2(n8264), .A(n8187), .ZN(n8182) );
  NAND2_X2 U8681 ( .A1(n8188), .A2(n8189), .ZN(n8187) );
  NAND2_X2 U8682 ( .A1(pipeline_regfile_data[478]), .A2(n6599), .ZN(n8189) );
  NAND2_X2 U8683 ( .A1(pipeline_regfile_data[414]), .A2(n8270), .ZN(n8188) );
  AND2_X1 U8684 ( .A1(n8190), .A2(n8191), .ZN(n8180) );
  AOI221_X2 U8685 ( .B1(pipeline_regfile_data[126]), .B2(n8249), .C1(
        pipeline_regfile_data[62]), .C2(n8251), .A(n8192), .ZN(n8191) );
  NAND2_X2 U8686 ( .A1(n8193), .A2(n8194), .ZN(n8192) );
  NAND2_X2 U8687 ( .A1(pipeline_regfile_data[254]), .A2(n8256), .ZN(n8194) );
  NAND2_X2 U8688 ( .A1(pipeline_regfile_data[190]), .A2(n8257), .ZN(n8193) );
  AOI221_X2 U8689 ( .B1(pipeline_regfile_data[94]), .B2(n8259), .C1(
        pipeline_regfile_data[30]), .C2(n8265), .A(n8195), .ZN(n8190) );
  NAND2_X2 U8690 ( .A1(n8196), .A2(n8197), .ZN(n8195) );
  NAND2_X2 U8691 ( .A1(pipeline_regfile_data[222]), .A2(n8268), .ZN(n8197) );
  NAND2_X2 U8692 ( .A1(pipeline_regfile_data[158]), .A2(n8270), .ZN(n8196) );
  AOI221_X2 U8693 ( .B1(pipeline_regfile_data[1022]), .B2(n6725), .C1(
        pipeline_regfile_data[766]), .C2(n6721), .A(n8198), .ZN(n8177) );
  INV_X4 U8694 ( .A(n8199), .ZN(n8198) );
  AOI221_X2 U8695 ( .B1(pipeline_regfile_data[574]), .B2(n6726), .C1(
        pipeline_regfile_data[830]), .C2(n6722), .A(n8200), .ZN(n8199) );
  AND2_X1 U8696 ( .A1(pipeline_regfile_data[638]), .A2(n6730), .ZN(n8200) );
  NAND2_X2 U8697 ( .A1(n8202), .A2(n8203), .ZN(n8201) );
  NAND2_X2 U8698 ( .A1(pipeline_regfile_data[670]), .A2(n6731), .ZN(n8203) );
  NAND2_X2 U8699 ( .A1(pipeline_regfile_data[894]), .A2(n6732), .ZN(n8202) );
  AOI221_X2 U8700 ( .B1(pipeline_regfile_data[542]), .B2(n6719), .C1(
        pipeline_regfile_data[990]), .C2(n6723), .A(n8204), .ZN(n8175) );
  INV_X4 U8701 ( .A(n8205), .ZN(n8204) );
  AOI221_X2 U8702 ( .B1(pipeline_regfile_data[798]), .B2(n6727), .C1(
        pipeline_regfile_data[606]), .C2(n6724), .A(n8206), .ZN(n8205) );
  AND2_X1 U8703 ( .A1(pipeline_regfile_data[862]), .A2(n6729), .ZN(n8206) );
  AOI221_X2 U8704 ( .B1(pipeline_regfile_data[959]), .B2(n6728), .C1(
        pipeline_regfile_data[703]), .C2(n6720), .A(n8211), .ZN(n8210) );
  OAI22_X2 U8705 ( .A1(n8212), .A2(n6695), .B1(n8213), .B2(n6663), .ZN(n8211)
         );
  AND2_X1 U8706 ( .A1(n8215), .A2(n8216), .ZN(n8213) );
  AOI221_X2 U8707 ( .B1(pipeline_regfile_data[383]), .B2(n8246), .C1(
        pipeline_regfile_data[319]), .C2(n8251), .A(n8217), .ZN(n8216) );
  NAND2_X2 U8708 ( .A1(n8218), .A2(n8219), .ZN(n8217) );
  NAND2_X2 U8709 ( .A1(pipeline_regfile_data[511]), .A2(n8255), .ZN(n8219) );
  NAND2_X2 U8710 ( .A1(pipeline_regfile_data[447]), .A2(n8257), .ZN(n8218) );
  AOI221_X2 U8711 ( .B1(pipeline_regfile_data[351]), .B2(n8258), .C1(
        pipeline_regfile_data[287]), .C2(n8264), .A(n8220), .ZN(n8215) );
  NAND2_X2 U8712 ( .A1(n8221), .A2(n8222), .ZN(n8220) );
  NAND2_X2 U8713 ( .A1(pipeline_regfile_data[479]), .A2(n6599), .ZN(n8222) );
  NAND2_X2 U8714 ( .A1(pipeline_regfile_data[415]), .A2(n8269), .ZN(n8221) );
  AND2_X1 U8715 ( .A1(n8224), .A2(n8225), .ZN(n8212) );
  AOI221_X2 U8716 ( .B1(pipeline_regfile_data[127]), .B2(n8246), .C1(
        pipeline_regfile_data[63]), .C2(n8251), .A(n8226), .ZN(n8225) );
  NAND2_X2 U8717 ( .A1(n8227), .A2(n8228), .ZN(n8226) );
  NAND2_X2 U8718 ( .A1(pipeline_regfile_data[255]), .A2(n8256), .ZN(n8228) );
  NAND2_X2 U8719 ( .A1(pipeline_regfile_data[191]), .A2(n8257), .ZN(n8227) );
  AOI221_X2 U8720 ( .B1(pipeline_regfile_data[95]), .B2(n8258), .C1(
        pipeline_regfile_data[31]), .C2(n8265), .A(n8229), .ZN(n8224) );
  NAND2_X2 U8721 ( .A1(n8230), .A2(n8231), .ZN(n8229) );
  NAND2_X2 U8722 ( .A1(pipeline_regfile_data[223]), .A2(n8268), .ZN(n8231) );
  NAND2_X2 U8723 ( .A1(pipeline_regfile_data[159]), .A2(n8269), .ZN(n8230) );
  AOI221_X2 U8724 ( .B1(pipeline_regfile_data[1023]), .B2(n6725), .C1(
        pipeline_regfile_data[767]), .C2(n6721), .A(n8233), .ZN(n8209) );
  INV_X4 U8725 ( .A(n8234), .ZN(n8233) );
  AOI221_X2 U8726 ( .B1(pipeline_regfile_data[575]), .B2(n6726), .C1(
        pipeline_regfile_data[831]), .C2(n6722), .A(n8235), .ZN(n8234) );
  AND2_X1 U8727 ( .A1(pipeline_regfile_data[639]), .A2(n6730), .ZN(n8235) );
  INV_X4 U8728 ( .A(n8236), .ZN(n7226) );
  NAND2_X2 U8729 ( .A1(n8238), .A2(n8239), .ZN(n8237) );
  NAND2_X2 U8730 ( .A1(pipeline_regfile_data[671]), .A2(n6731), .ZN(n8239) );
  NAND2_X2 U8731 ( .A1(pipeline_regfile_data[895]), .A2(n6732), .ZN(n8238) );
  AOI221_X2 U8732 ( .B1(pipeline_regfile_data[543]), .B2(n6719), .C1(
        pipeline_regfile_data[991]), .C2(n6723), .A(n8241), .ZN(n8207) );
  INV_X4 U8733 ( .A(n8242), .ZN(n8241) );
  AOI221_X2 U8734 ( .B1(pipeline_regfile_data[799]), .B2(n6727), .C1(
        pipeline_regfile_data[607]), .C2(n6724), .A(n8243), .ZN(n8242) );
  AND2_X1 U8735 ( .A1(pipeline_regfile_data[863]), .A2(n6729), .ZN(n8243) );
  NAND3_X1 U8736 ( .A1(pipeline_regfile_N17), .A2(n702), .A3(n9658), .ZN(n8236) );
  AOI221_X2 U8737 ( .B1(pipeline_regfile_data[928]), .B2(n6767), .C1(
        pipeline_regfile_data[672]), .C2(n6764), .A(n8276), .ZN(n8275) );
  OAI22_X2 U8738 ( .A1(n8277), .A2(n8278), .B1(n8279), .B2(n9306), .ZN(n8276)
         );
  AND2_X1 U8739 ( .A1(n8280), .A2(n8281), .ZN(n8279) );
  AOI221_X2 U8740 ( .B1(pipeline_regfile_data[352]), .B2(n9310), .C1(
        pipeline_regfile_data[288]), .C2(n9316), .A(n8282), .ZN(n8281) );
  NAND2_X2 U8741 ( .A1(n8283), .A2(n8284), .ZN(n8282) );
  NAND2_X2 U8742 ( .A1(pipeline_regfile_data[480]), .A2(n9318), .ZN(n8284) );
  NAND2_X2 U8743 ( .A1(pipeline_regfile_data[416]), .A2(n9321), .ZN(n8283) );
  AOI221_X2 U8744 ( .B1(pipeline_regfile_data[320]), .B2(n9325), .C1(
        pipeline_regfile_data[256]), .C2(n9327), .A(n8286), .ZN(n8280) );
  NAND2_X2 U8745 ( .A1(n8287), .A2(n8288), .ZN(n8286) );
  NAND2_X2 U8746 ( .A1(pipeline_regfile_data[448]), .A2(n9328), .ZN(n8288) );
  NAND2_X2 U8747 ( .A1(pipeline_regfile_data[384]), .A2(n9330), .ZN(n8287) );
  AND2_X1 U8748 ( .A1(n8289), .A2(n8290), .ZN(n8277) );
  AOI221_X2 U8749 ( .B1(pipeline_regfile_data[96]), .B2(n9310), .C1(
        pipeline_regfile_data[32]), .C2(n9316), .A(n8291), .ZN(n8290) );
  NAND2_X2 U8750 ( .A1(n8292), .A2(n8293), .ZN(n8291) );
  NAND2_X2 U8751 ( .A1(pipeline_regfile_data[224]), .A2(n9318), .ZN(n8293) );
  NAND2_X2 U8752 ( .A1(pipeline_regfile_data[160]), .A2(n9321), .ZN(n8292) );
  AOI221_X2 U8753 ( .B1(pipeline_regfile_data[64]), .B2(n9325), .C1(
        pipeline_regfile_data[0]), .C2(n9326), .A(n8294), .ZN(n8289) );
  NAND2_X2 U8754 ( .A1(n8295), .A2(n8296), .ZN(n8294) );
  NAND2_X2 U8755 ( .A1(pipeline_regfile_data[192]), .A2(n9328), .ZN(n8296) );
  NAND2_X2 U8756 ( .A1(pipeline_regfile_data[128]), .A2(n9330), .ZN(n8295) );
  AOI221_X2 U8757 ( .B1(pipeline_regfile_data[992]), .B2(n6765), .C1(
        pipeline_regfile_data[736]), .C2(n6761), .A(n8297), .ZN(n8274) );
  INV_X4 U8758 ( .A(n8298), .ZN(n8297) );
  AOI221_X2 U8759 ( .B1(pipeline_regfile_data[544]), .B2(n8299), .C1(
        pipeline_regfile_data[800]), .C2(n8300), .A(n8301), .ZN(n8298) );
  AND2_X1 U8760 ( .A1(pipeline_regfile_data[608]), .A2(n8302), .ZN(n8301) );
  NAND2_X2 U8761 ( .A1(n8304), .A2(n8305), .ZN(n8303) );
  NAND2_X2 U8762 ( .A1(pipeline_regfile_data[640]), .A2(n6769), .ZN(n8305) );
  NAND2_X2 U8763 ( .A1(pipeline_regfile_data[864]), .A2(n6770), .ZN(n8304) );
  AOI221_X2 U8764 ( .B1(pipeline_regfile_data[512]), .B2(n6709), .C1(
        pipeline_regfile_data[960]), .C2(n6763), .A(n8306), .ZN(n8272) );
  INV_X4 U8765 ( .A(n8307), .ZN(n8306) );
  AOI221_X2 U8766 ( .B1(pipeline_regfile_data[768]), .B2(n6766), .C1(
        pipeline_regfile_data[576]), .C2(n6762), .A(n8308), .ZN(n8307) );
  AND2_X1 U8767 ( .A1(pipeline_regfile_data[832]), .A2(n6768), .ZN(n8308) );
  OAI22_X2 U8768 ( .A1(n8313), .A2(n8278), .B1(n8314), .B2(n9306), .ZN(n8312)
         );
  AOI221_X2 U8769 ( .B1(pipeline_regfile_data[353]), .B2(n9310), .C1(
        pipeline_regfile_data[289]), .C2(n9316), .A(n8317), .ZN(n8316) );
  NAND2_X2 U8770 ( .A1(n8318), .A2(n8319), .ZN(n8317) );
  NAND2_X2 U8771 ( .A1(pipeline_regfile_data[481]), .A2(n9318), .ZN(n8319) );
  NAND2_X2 U8772 ( .A1(pipeline_regfile_data[417]), .A2(n9321), .ZN(n8318) );
  AOI221_X2 U8773 ( .B1(pipeline_regfile_data[321]), .B2(n9325), .C1(
        pipeline_regfile_data[257]), .C2(n9326), .A(n8320), .ZN(n8315) );
  NAND2_X2 U8774 ( .A1(n8321), .A2(n8322), .ZN(n8320) );
  NAND2_X2 U8775 ( .A1(pipeline_regfile_data[449]), .A2(n9328), .ZN(n8322) );
  NAND2_X2 U8776 ( .A1(pipeline_regfile_data[385]), .A2(n7171), .ZN(n8321) );
  AND2_X1 U8777 ( .A1(n8323), .A2(n8324), .ZN(n8313) );
  AOI221_X2 U8778 ( .B1(pipeline_regfile_data[97]), .B2(n9310), .C1(
        pipeline_regfile_data[33]), .C2(n9316), .A(n8325), .ZN(n8324) );
  NAND2_X2 U8779 ( .A1(n8326), .A2(n8327), .ZN(n8325) );
  NAND2_X2 U8780 ( .A1(pipeline_regfile_data[225]), .A2(n9318), .ZN(n8327) );
  NAND2_X2 U8781 ( .A1(pipeline_regfile_data[161]), .A2(n9321), .ZN(n8326) );
  AOI221_X2 U8782 ( .B1(pipeline_regfile_data[65]), .B2(n9325), .C1(
        pipeline_regfile_data[1]), .C2(n9326), .A(n8328), .ZN(n8323) );
  NAND2_X2 U8783 ( .A1(n8329), .A2(n8330), .ZN(n8328) );
  NAND2_X2 U8784 ( .A1(pipeline_regfile_data[193]), .A2(n9328), .ZN(n8330) );
  NAND2_X2 U8785 ( .A1(pipeline_regfile_data[129]), .A2(n7171), .ZN(n8329) );
  AOI221_X2 U8786 ( .B1(pipeline_regfile_data[993]), .B2(n6765), .C1(
        pipeline_regfile_data[737]), .C2(n6761), .A(n8331), .ZN(n8311) );
  INV_X4 U8787 ( .A(n8332), .ZN(n8331) );
  AOI221_X2 U8788 ( .B1(pipeline_regfile_data[545]), .B2(n8299), .C1(
        pipeline_regfile_data[801]), .C2(n8300), .A(n8333), .ZN(n8332) );
  AND2_X1 U8789 ( .A1(pipeline_regfile_data[609]), .A2(n8302), .ZN(n8333) );
  AOI221_X2 U8790 ( .B1(pipeline_regfile_data[705]), .B2(n6773), .C1(
        pipeline_regfile_data[897]), .C2(n6772), .A(n8334), .ZN(n8310) );
  NAND2_X2 U8791 ( .A1(n8335), .A2(n8336), .ZN(n8334) );
  NAND2_X2 U8792 ( .A1(pipeline_regfile_data[641]), .A2(n6769), .ZN(n8336) );
  NAND2_X2 U8793 ( .A1(pipeline_regfile_data[865]), .A2(n6770), .ZN(n8335) );
  AOI221_X2 U8794 ( .B1(pipeline_regfile_data[513]), .B2(n6709), .C1(
        pipeline_regfile_data[961]), .C2(n6763), .A(n8337), .ZN(n8309) );
  INV_X4 U8795 ( .A(n8338), .ZN(n8337) );
  AOI221_X2 U8796 ( .B1(pipeline_regfile_data[769]), .B2(n6766), .C1(
        pipeline_regfile_data[577]), .C2(n6762), .A(n8339), .ZN(n8338) );
  AND2_X1 U8797 ( .A1(pipeline_regfile_data[833]), .A2(n6768), .ZN(n8339) );
  AOI221_X2 U8798 ( .B1(pipeline_regfile_data[930]), .B2(n6767), .C1(
        pipeline_regfile_data[674]), .C2(n6764), .A(n8344), .ZN(n8343) );
  OAI22_X2 U8799 ( .A1(n8345), .A2(n8278), .B1(n8346), .B2(n9306), .ZN(n8344)
         );
  AND2_X1 U8800 ( .A1(n8347), .A2(n8348), .ZN(n8346) );
  AOI221_X2 U8801 ( .B1(pipeline_regfile_data[354]), .B2(n9310), .C1(
        pipeline_regfile_data[290]), .C2(n9316), .A(n8349), .ZN(n8348) );
  NAND2_X2 U8802 ( .A1(n8350), .A2(n8351), .ZN(n8349) );
  NAND2_X2 U8803 ( .A1(pipeline_regfile_data[482]), .A2(n9318), .ZN(n8351) );
  NAND2_X2 U8804 ( .A1(pipeline_regfile_data[418]), .A2(n9321), .ZN(n8350) );
  AOI221_X2 U8805 ( .B1(pipeline_regfile_data[322]), .B2(n9325), .C1(
        pipeline_regfile_data[258]), .C2(n9326), .A(n8352), .ZN(n8347) );
  NAND2_X2 U8806 ( .A1(n8353), .A2(n8354), .ZN(n8352) );
  NAND2_X2 U8807 ( .A1(pipeline_regfile_data[450]), .A2(n9328), .ZN(n8354) );
  NAND2_X2 U8808 ( .A1(pipeline_regfile_data[386]), .A2(n7171), .ZN(n8353) );
  AND2_X1 U8809 ( .A1(n8355), .A2(n8356), .ZN(n8345) );
  AOI221_X2 U8810 ( .B1(pipeline_regfile_data[98]), .B2(n9310), .C1(
        pipeline_regfile_data[34]), .C2(n9316), .A(n8357), .ZN(n8356) );
  NAND2_X2 U8811 ( .A1(n8358), .A2(n8359), .ZN(n8357) );
  NAND2_X2 U8812 ( .A1(pipeline_regfile_data[226]), .A2(n9318), .ZN(n8359) );
  NAND2_X2 U8813 ( .A1(pipeline_regfile_data[162]), .A2(n9321), .ZN(n8358) );
  AOI221_X2 U8814 ( .B1(pipeline_regfile_data[66]), .B2(n9325), .C1(
        pipeline_regfile_data[2]), .C2(n9326), .A(n8360), .ZN(n8355) );
  NAND2_X2 U8815 ( .A1(n8361), .A2(n8362), .ZN(n8360) );
  NAND2_X2 U8816 ( .A1(pipeline_regfile_data[194]), .A2(n9328), .ZN(n8362) );
  NAND2_X2 U8817 ( .A1(pipeline_regfile_data[130]), .A2(n7171), .ZN(n8361) );
  AOI221_X2 U8818 ( .B1(pipeline_regfile_data[994]), .B2(n6765), .C1(
        pipeline_regfile_data[738]), .C2(n6761), .A(n8363), .ZN(n8342) );
  INV_X4 U8819 ( .A(n8364), .ZN(n8363) );
  AOI221_X2 U8820 ( .B1(pipeline_regfile_data[546]), .B2(n8299), .C1(
        pipeline_regfile_data[802]), .C2(n8300), .A(n8365), .ZN(n8364) );
  AND2_X1 U8821 ( .A1(pipeline_regfile_data[610]), .A2(n8302), .ZN(n8365) );
  AOI221_X2 U8822 ( .B1(pipeline_regfile_data[706]), .B2(n6773), .C1(
        pipeline_regfile_data[898]), .C2(n6772), .A(n8366), .ZN(n8341) );
  NAND2_X2 U8823 ( .A1(n8367), .A2(n8368), .ZN(n8366) );
  NAND2_X2 U8824 ( .A1(pipeline_regfile_data[642]), .A2(n6769), .ZN(n8368) );
  NAND2_X2 U8825 ( .A1(pipeline_regfile_data[866]), .A2(n6770), .ZN(n8367) );
  AOI221_X2 U8826 ( .B1(pipeline_regfile_data[514]), .B2(n6709), .C1(
        pipeline_regfile_data[962]), .C2(n6763), .A(n8369), .ZN(n8340) );
  INV_X4 U8827 ( .A(n8370), .ZN(n8369) );
  AOI221_X2 U8828 ( .B1(pipeline_regfile_data[770]), .B2(n6766), .C1(
        pipeline_regfile_data[578]), .C2(n6762), .A(n8371), .ZN(n8370) );
  AND2_X1 U8829 ( .A1(pipeline_regfile_data[834]), .A2(n6768), .ZN(n8371) );
  OAI22_X2 U8830 ( .A1(n8377), .A2(n9305), .B1(n8378), .B2(n9306), .ZN(n8376)
         );
  AOI221_X2 U8831 ( .B1(pipeline_regfile_data[355]), .B2(n9310), .C1(
        pipeline_regfile_data[291]), .C2(n9316), .A(n8381), .ZN(n8380) );
  NAND2_X2 U8832 ( .A1(n8382), .A2(n8383), .ZN(n8381) );
  NAND2_X2 U8833 ( .A1(pipeline_regfile_data[483]), .A2(n9318), .ZN(n8383) );
  NAND2_X2 U8834 ( .A1(pipeline_regfile_data[419]), .A2(n9321), .ZN(n8382) );
  AOI221_X2 U8835 ( .B1(pipeline_regfile_data[323]), .B2(n9325), .C1(
        pipeline_regfile_data[259]), .C2(n9326), .A(n8384), .ZN(n8379) );
  NAND2_X2 U8836 ( .A1(n8385), .A2(n8386), .ZN(n8384) );
  NAND2_X2 U8837 ( .A1(pipeline_regfile_data[451]), .A2(n9328), .ZN(n8386) );
  NAND2_X2 U8838 ( .A1(pipeline_regfile_data[387]), .A2(n9329), .ZN(n8385) );
  AND2_X1 U8839 ( .A1(n8387), .A2(n8388), .ZN(n8377) );
  AOI221_X2 U8840 ( .B1(pipeline_regfile_data[99]), .B2(n9310), .C1(
        pipeline_regfile_data[35]), .C2(n9316), .A(n8389), .ZN(n8388) );
  NAND2_X2 U8841 ( .A1(n8390), .A2(n8391), .ZN(n8389) );
  NAND2_X2 U8842 ( .A1(pipeline_regfile_data[227]), .A2(n9318), .ZN(n8391) );
  NAND2_X2 U8843 ( .A1(pipeline_regfile_data[163]), .A2(n9321), .ZN(n8390) );
  AOI221_X2 U8844 ( .B1(pipeline_regfile_data[67]), .B2(n9325), .C1(
        pipeline_regfile_data[3]), .C2(n9326), .A(n8392), .ZN(n8387) );
  NAND2_X2 U8845 ( .A1(n8393), .A2(n8394), .ZN(n8392) );
  NAND2_X2 U8846 ( .A1(pipeline_regfile_data[195]), .A2(n9328), .ZN(n8394) );
  NAND2_X2 U8847 ( .A1(pipeline_regfile_data[131]), .A2(n9330), .ZN(n8393) );
  AOI221_X2 U8848 ( .B1(pipeline_regfile_data[995]), .B2(n6765), .C1(
        pipeline_regfile_data[739]), .C2(n6761), .A(n6933), .ZN(n8374) );
  AOI221_X2 U8849 ( .B1(pipeline_regfile_data[707]), .B2(n6773), .C1(
        pipeline_regfile_data[899]), .C2(n6772), .A(n8395), .ZN(n8373) );
  NAND2_X2 U8850 ( .A1(n8396), .A2(n8397), .ZN(n8395) );
  NAND2_X2 U8851 ( .A1(pipeline_regfile_data[643]), .A2(n6769), .ZN(n8397) );
  NAND2_X2 U8852 ( .A1(pipeline_regfile_data[867]), .A2(n6770), .ZN(n8396) );
  AOI221_X2 U8853 ( .B1(pipeline_regfile_data[515]), .B2(n6709), .C1(
        pipeline_regfile_data[963]), .C2(n6763), .A(n8398), .ZN(n8372) );
  INV_X4 U8854 ( .A(n8399), .ZN(n8398) );
  AOI221_X2 U8855 ( .B1(pipeline_regfile_data[771]), .B2(n6766), .C1(
        pipeline_regfile_data[579]), .C2(n6762), .A(n8400), .ZN(n8399) );
  AND2_X1 U8856 ( .A1(pipeline_regfile_data[835]), .A2(n6768), .ZN(n8400) );
  AOI221_X2 U8857 ( .B1(pipeline_regfile_data[356]), .B2(n9310), .C1(
        pipeline_regfile_data[292]), .C2(n9316), .A(n8410), .ZN(n8409) );
  NAND2_X2 U8858 ( .A1(n8411), .A2(n8412), .ZN(n8410) );
  NAND2_X2 U8859 ( .A1(pipeline_regfile_data[484]), .A2(n9320), .ZN(n8412) );
  NAND2_X2 U8860 ( .A1(pipeline_regfile_data[420]), .A2(n9321), .ZN(n8411) );
  AOI221_X2 U8861 ( .B1(pipeline_regfile_data[324]), .B2(n9325), .C1(
        pipeline_regfile_data[260]), .C2(n9326), .A(n8413), .ZN(n8408) );
  NAND2_X2 U8862 ( .A1(n8414), .A2(n8415), .ZN(n8413) );
  NAND2_X2 U8863 ( .A1(pipeline_regfile_data[452]), .A2(n9328), .ZN(n8415) );
  NAND2_X2 U8864 ( .A1(pipeline_regfile_data[388]), .A2(n9330), .ZN(n8414) );
  AOI221_X2 U8865 ( .B1(pipeline_regfile_data[100]), .B2(n9310), .C1(
        pipeline_regfile_data[36]), .C2(n9316), .A(n8418), .ZN(n8417) );
  NAND2_X2 U8866 ( .A1(n8419), .A2(n8420), .ZN(n8418) );
  NAND2_X2 U8867 ( .A1(pipeline_regfile_data[228]), .A2(n9320), .ZN(n8420) );
  NAND2_X2 U8868 ( .A1(pipeline_regfile_data[164]), .A2(n9321), .ZN(n8419) );
  AOI221_X2 U8869 ( .B1(pipeline_regfile_data[68]), .B2(n9325), .C1(
        pipeline_regfile_data[4]), .C2(n9326), .A(n8421), .ZN(n8416) );
  NAND2_X2 U8870 ( .A1(n8422), .A2(n8423), .ZN(n8421) );
  NAND2_X2 U8871 ( .A1(pipeline_regfile_data[196]), .A2(n9328), .ZN(n8423) );
  NAND2_X2 U8872 ( .A1(pipeline_regfile_data[132]), .A2(n9330), .ZN(n8422) );
  AOI221_X2 U8873 ( .B1(pipeline_regfile_data[996]), .B2(n6765), .C1(
        pipeline_regfile_data[740]), .C2(n6761), .A(n8424), .ZN(n8403) );
  AOI221_X2 U8874 ( .B1(pipeline_regfile_data[548]), .B2(n8299), .C1(
        pipeline_regfile_data[804]), .C2(n8300), .A(n8426), .ZN(n8425) );
  AOI221_X2 U8875 ( .B1(pipeline_regfile_data[708]), .B2(n6773), .C1(
        pipeline_regfile_data[900]), .C2(n6772), .A(n8427), .ZN(n8402) );
  NAND2_X2 U8876 ( .A1(n8428), .A2(n8429), .ZN(n8427) );
  NAND2_X2 U8877 ( .A1(pipeline_regfile_data[644]), .A2(n6769), .ZN(n8429) );
  NAND2_X2 U8878 ( .A1(pipeline_regfile_data[868]), .A2(n6770), .ZN(n8428) );
  AOI221_X2 U8879 ( .B1(pipeline_regfile_data[516]), .B2(n6709), .C1(
        pipeline_regfile_data[964]), .C2(n6763), .A(n8430), .ZN(n8401) );
  AOI221_X2 U8880 ( .B1(pipeline_regfile_data[772]), .B2(n6766), .C1(
        pipeline_regfile_data[580]), .C2(n6762), .A(n8432), .ZN(n8431) );
  AND2_X1 U8881 ( .A1(pipeline_regfile_data[836]), .A2(n6768), .ZN(n8432) );
  AOI221_X2 U8882 ( .B1(pipeline_regfile_data[933]), .B2(n6767), .C1(
        pipeline_regfile_data[677]), .C2(n6764), .A(n8437), .ZN(n8436) );
  OAI22_X2 U8883 ( .A1(n8438), .A2(n8278), .B1(n8439), .B2(n9306), .ZN(n8437)
         );
  AND2_X1 U8884 ( .A1(n8440), .A2(n8441), .ZN(n8439) );
  AOI221_X2 U8885 ( .B1(pipeline_regfile_data[357]), .B2(n9310), .C1(
        pipeline_regfile_data[293]), .C2(n9316), .A(n8442), .ZN(n8441) );
  NAND2_X2 U8886 ( .A1(n8443), .A2(n8444), .ZN(n8442) );
  NAND2_X2 U8887 ( .A1(pipeline_regfile_data[485]), .A2(n9318), .ZN(n8444) );
  NAND2_X2 U8888 ( .A1(pipeline_regfile_data[421]), .A2(n9321), .ZN(n8443) );
  AOI221_X2 U8889 ( .B1(pipeline_regfile_data[325]), .B2(n9325), .C1(
        pipeline_regfile_data[261]), .C2(n9326), .A(n8445), .ZN(n8440) );
  NAND2_X2 U8890 ( .A1(pipeline_regfile_data[453]), .A2(n9328), .ZN(n8447) );
  NAND2_X2 U8891 ( .A1(pipeline_regfile_data[389]), .A2(n9330), .ZN(n8446) );
  AND2_X1 U8892 ( .A1(n8448), .A2(n8449), .ZN(n8438) );
  AOI221_X2 U8893 ( .B1(pipeline_regfile_data[101]), .B2(n9310), .C1(
        pipeline_regfile_data[37]), .C2(n9316), .A(n8450), .ZN(n8449) );
  NAND2_X2 U8894 ( .A1(n8451), .A2(n8452), .ZN(n8450) );
  NAND2_X2 U8895 ( .A1(pipeline_regfile_data[229]), .A2(n9318), .ZN(n8452) );
  NAND2_X2 U8896 ( .A1(pipeline_regfile_data[165]), .A2(n9321), .ZN(n8451) );
  AOI221_X2 U8897 ( .B1(pipeline_regfile_data[69]), .B2(n9325), .C1(
        pipeline_regfile_data[5]), .C2(n9326), .A(n8453), .ZN(n8448) );
  NAND2_X2 U8898 ( .A1(n8454), .A2(n8455), .ZN(n8453) );
  NAND2_X2 U8899 ( .A1(pipeline_regfile_data[197]), .A2(n9328), .ZN(n8455) );
  NAND2_X2 U8900 ( .A1(pipeline_regfile_data[133]), .A2(n9329), .ZN(n8454) );
  AOI221_X2 U8901 ( .B1(pipeline_regfile_data[997]), .B2(n6765), .C1(
        pipeline_regfile_data[741]), .C2(n6761), .A(n8456), .ZN(n8435) );
  INV_X4 U8902 ( .A(n8457), .ZN(n8456) );
  AOI221_X2 U8903 ( .B1(pipeline_regfile_data[549]), .B2(n8299), .C1(
        pipeline_regfile_data[805]), .C2(n8300), .A(n8458), .ZN(n8457) );
  AND2_X1 U8904 ( .A1(pipeline_regfile_data[613]), .A2(n8302), .ZN(n8458) );
  NAND2_X2 U8905 ( .A1(n8460), .A2(n8461), .ZN(n8459) );
  NAND2_X2 U8906 ( .A1(pipeline_regfile_data[645]), .A2(n6769), .ZN(n8461) );
  NAND2_X2 U8907 ( .A1(pipeline_regfile_data[869]), .A2(n6770), .ZN(n8460) );
  AOI221_X2 U8908 ( .B1(pipeline_regfile_data[517]), .B2(n6709), .C1(
        pipeline_regfile_data[965]), .C2(n6763), .A(n8462), .ZN(n8433) );
  INV_X4 U8909 ( .A(n8463), .ZN(n8462) );
  AOI221_X2 U8910 ( .B1(pipeline_regfile_data[773]), .B2(n6766), .C1(
        pipeline_regfile_data[581]), .C2(n6762), .A(n8464), .ZN(n8463) );
  AND2_X1 U8911 ( .A1(pipeline_regfile_data[837]), .A2(n6768), .ZN(n8464) );
  AOI221_X2 U8912 ( .B1(pipeline_regfile_data[934]), .B2(n6767), .C1(
        pipeline_regfile_data[678]), .C2(n6764), .A(n8469), .ZN(n8468) );
  OAI22_X2 U8913 ( .A1(n8470), .A2(n8278), .B1(n8471), .B2(n9306), .ZN(n8469)
         );
  AND2_X1 U8914 ( .A1(n8472), .A2(n8473), .ZN(n8471) );
  AOI221_X2 U8915 ( .B1(pipeline_regfile_data[358]), .B2(n9310), .C1(
        pipeline_regfile_data[294]), .C2(n9316), .A(n8474), .ZN(n8473) );
  NAND2_X2 U8916 ( .A1(n8475), .A2(n8476), .ZN(n8474) );
  NAND2_X2 U8917 ( .A1(pipeline_regfile_data[486]), .A2(n9318), .ZN(n8476) );
  NAND2_X2 U8918 ( .A1(pipeline_regfile_data[422]), .A2(n9321), .ZN(n8475) );
  AOI221_X2 U8919 ( .B1(pipeline_regfile_data[326]), .B2(n9325), .C1(
        pipeline_regfile_data[262]), .C2(n9327), .A(n8477), .ZN(n8472) );
  NAND2_X2 U8920 ( .A1(n8478), .A2(n8479), .ZN(n8477) );
  NAND2_X2 U8921 ( .A1(pipeline_regfile_data[454]), .A2(n9328), .ZN(n8479) );
  NAND2_X2 U8922 ( .A1(pipeline_regfile_data[390]), .A2(n7171), .ZN(n8478) );
  AND2_X1 U8923 ( .A1(n8480), .A2(n8481), .ZN(n8470) );
  AOI221_X2 U8924 ( .B1(pipeline_regfile_data[102]), .B2(n9309), .C1(
        pipeline_regfile_data[38]), .C2(n9315), .A(n8482), .ZN(n8481) );
  NAND2_X2 U8925 ( .A1(n8483), .A2(n8484), .ZN(n8482) );
  NAND2_X2 U8926 ( .A1(pipeline_regfile_data[230]), .A2(n9318), .ZN(n8484) );
  NAND2_X2 U8927 ( .A1(pipeline_regfile_data[166]), .A2(n9321), .ZN(n8483) );
  AOI221_X2 U8928 ( .B1(pipeline_regfile_data[70]), .B2(n9324), .C1(
        pipeline_regfile_data[6]), .C2(n9327), .A(n8485), .ZN(n8480) );
  NAND2_X2 U8929 ( .A1(n8486), .A2(n8487), .ZN(n8485) );
  NAND2_X2 U8930 ( .A1(pipeline_regfile_data[198]), .A2(n9328), .ZN(n8487) );
  NAND2_X2 U8931 ( .A1(pipeline_regfile_data[134]), .A2(n7171), .ZN(n8486) );
  AOI221_X2 U8932 ( .B1(pipeline_regfile_data[998]), .B2(n6765), .C1(
        pipeline_regfile_data[742]), .C2(n6761), .A(n8488), .ZN(n8467) );
  INV_X4 U8933 ( .A(n8489), .ZN(n8488) );
  AOI221_X2 U8934 ( .B1(pipeline_regfile_data[550]), .B2(n8299), .C1(
        pipeline_regfile_data[806]), .C2(n8300), .A(n8490), .ZN(n8489) );
  AND2_X1 U8935 ( .A1(pipeline_regfile_data[614]), .A2(n8302), .ZN(n8490) );
  AOI221_X2 U8936 ( .B1(pipeline_regfile_data[710]), .B2(n6773), .C1(
        pipeline_regfile_data[902]), .C2(n6772), .A(n8491), .ZN(n8466) );
  NAND2_X2 U8937 ( .A1(n8492), .A2(n8493), .ZN(n8491) );
  NAND2_X2 U8938 ( .A1(pipeline_regfile_data[646]), .A2(n6769), .ZN(n8493) );
  NAND2_X2 U8939 ( .A1(pipeline_regfile_data[870]), .A2(n6770), .ZN(n8492) );
  AOI221_X2 U8940 ( .B1(pipeline_regfile_data[518]), .B2(n6709), .C1(
        pipeline_regfile_data[966]), .C2(n6763), .A(n8494), .ZN(n8465) );
  INV_X4 U8941 ( .A(n8495), .ZN(n8494) );
  AOI221_X2 U8942 ( .B1(pipeline_regfile_data[774]), .B2(n6766), .C1(
        pipeline_regfile_data[582]), .C2(n6762), .A(n8496), .ZN(n8495) );
  AND2_X1 U8943 ( .A1(pipeline_regfile_data[838]), .A2(n6768), .ZN(n8496) );
  AOI221_X2 U8944 ( .B1(pipeline_regfile_data[935]), .B2(n6767), .C1(
        pipeline_regfile_data[679]), .C2(n6764), .A(n8501), .ZN(n8500) );
  AND2_X1 U8945 ( .A1(n8504), .A2(n8505), .ZN(n8503) );
  AOI221_X2 U8946 ( .B1(pipeline_regfile_data[359]), .B2(n9309), .C1(
        pipeline_regfile_data[295]), .C2(n9315), .A(n8506), .ZN(n8505) );
  NAND2_X2 U8947 ( .A1(n8507), .A2(n8508), .ZN(n8506) );
  NAND2_X2 U8948 ( .A1(pipeline_regfile_data[487]), .A2(n9318), .ZN(n8508) );
  NAND2_X2 U8949 ( .A1(pipeline_regfile_data[423]), .A2(n9321), .ZN(n8507) );
  AOI221_X2 U8950 ( .B1(pipeline_regfile_data[327]), .B2(n9324), .C1(
        pipeline_regfile_data[263]), .C2(n9327), .A(n8509), .ZN(n8504) );
  NAND2_X2 U8951 ( .A1(n8510), .A2(n8511), .ZN(n8509) );
  NAND2_X2 U8952 ( .A1(pipeline_regfile_data[455]), .A2(n9328), .ZN(n8511) );
  NAND2_X2 U8953 ( .A1(pipeline_regfile_data[391]), .A2(n7171), .ZN(n8510) );
  AND2_X1 U8954 ( .A1(n8512), .A2(n8513), .ZN(n8502) );
  AOI221_X2 U8955 ( .B1(pipeline_regfile_data[103]), .B2(n9308), .C1(
        pipeline_regfile_data[39]), .C2(n9315), .A(n8514), .ZN(n8513) );
  NAND2_X2 U8956 ( .A1(n8515), .A2(n8516), .ZN(n8514) );
  NAND2_X2 U8957 ( .A1(pipeline_regfile_data[231]), .A2(n9318), .ZN(n8516) );
  NAND2_X2 U8958 ( .A1(pipeline_regfile_data[167]), .A2(n9321), .ZN(n8515) );
  AOI221_X2 U8959 ( .B1(pipeline_regfile_data[71]), .B2(n9324), .C1(
        pipeline_regfile_data[7]), .C2(n9327), .A(n8517), .ZN(n8512) );
  NAND2_X2 U8960 ( .A1(n8518), .A2(n8519), .ZN(n8517) );
  NAND2_X2 U8961 ( .A1(pipeline_regfile_data[199]), .A2(n9328), .ZN(n8519) );
  NAND2_X2 U8962 ( .A1(pipeline_regfile_data[135]), .A2(n9330), .ZN(n8518) );
  AOI221_X2 U8963 ( .B1(pipeline_regfile_data[999]), .B2(n6765), .C1(
        pipeline_regfile_data[743]), .C2(n6761), .A(n8520), .ZN(n8499) );
  INV_X4 U8964 ( .A(n8521), .ZN(n8520) );
  AOI221_X2 U8965 ( .B1(pipeline_regfile_data[551]), .B2(n8299), .C1(
        pipeline_regfile_data[807]), .C2(n8300), .A(n8522), .ZN(n8521) );
  AND2_X1 U8966 ( .A1(pipeline_regfile_data[615]), .A2(n8302), .ZN(n8522) );
  AOI221_X2 U8967 ( .B1(pipeline_regfile_data[711]), .B2(n6773), .C1(
        pipeline_regfile_data[903]), .C2(n6772), .A(n8523), .ZN(n8498) );
  NAND2_X2 U8968 ( .A1(n8524), .A2(n8525), .ZN(n8523) );
  NAND2_X2 U8969 ( .A1(pipeline_regfile_data[647]), .A2(n6769), .ZN(n8525) );
  NAND2_X2 U8970 ( .A1(pipeline_regfile_data[871]), .A2(n6770), .ZN(n8524) );
  AOI221_X2 U8971 ( .B1(pipeline_regfile_data[519]), .B2(n6709), .C1(
        pipeline_regfile_data[967]), .C2(n6763), .A(n8526), .ZN(n8497) );
  INV_X4 U8972 ( .A(n8527), .ZN(n8526) );
  AOI221_X2 U8973 ( .B1(pipeline_regfile_data[775]), .B2(n6766), .C1(
        pipeline_regfile_data[583]), .C2(n6762), .A(n8528), .ZN(n8527) );
  AND2_X1 U8974 ( .A1(pipeline_regfile_data[839]), .A2(n6768), .ZN(n8528) );
  AOI221_X2 U8975 ( .B1(pipeline_regfile_data[936]), .B2(n6767), .C1(
        pipeline_regfile_data[680]), .C2(n6764), .A(n8533), .ZN(n8532) );
  OAI22_X2 U8976 ( .A1(n8534), .A2(n8278), .B1(n8535), .B2(n9306), .ZN(n8533)
         );
  AND2_X1 U8977 ( .A1(n8536), .A2(n8537), .ZN(n8535) );
  AOI221_X2 U8978 ( .B1(pipeline_regfile_data[360]), .B2(n9308), .C1(
        pipeline_regfile_data[296]), .C2(n9315), .A(n8538), .ZN(n8537) );
  NAND2_X2 U8979 ( .A1(n8539), .A2(n8540), .ZN(n8538) );
  NAND2_X2 U8980 ( .A1(pipeline_regfile_data[488]), .A2(n9318), .ZN(n8540) );
  NAND2_X2 U8981 ( .A1(pipeline_regfile_data[424]), .A2(n9321), .ZN(n8539) );
  NAND2_X2 U8982 ( .A1(n8542), .A2(n8543), .ZN(n8541) );
  NAND2_X2 U8983 ( .A1(pipeline_regfile_data[456]), .A2(n9328), .ZN(n8543) );
  NAND2_X2 U8984 ( .A1(pipeline_regfile_data[392]), .A2(n9332), .ZN(n8542) );
  AND2_X1 U8985 ( .A1(n8544), .A2(n8545), .ZN(n8534) );
  AOI221_X2 U8986 ( .B1(pipeline_regfile_data[104]), .B2(n9309), .C1(
        pipeline_regfile_data[40]), .C2(n9315), .A(n8546), .ZN(n8545) );
  NAND2_X2 U8987 ( .A1(n8547), .A2(n8548), .ZN(n8546) );
  NAND2_X2 U8988 ( .A1(pipeline_regfile_data[232]), .A2(n9318), .ZN(n8548) );
  NAND2_X2 U8989 ( .A1(pipeline_regfile_data[168]), .A2(n9321), .ZN(n8547) );
  AOI221_X2 U8990 ( .B1(pipeline_regfile_data[72]), .B2(n9324), .C1(
        pipeline_regfile_data[8]), .C2(n9327), .A(n8549), .ZN(n8544) );
  NAND2_X2 U8991 ( .A1(n8550), .A2(n8551), .ZN(n8549) );
  NAND2_X2 U8992 ( .A1(pipeline_regfile_data[200]), .A2(n9328), .ZN(n8551) );
  NAND2_X2 U8993 ( .A1(pipeline_regfile_data[136]), .A2(n9330), .ZN(n8550) );
  AOI221_X2 U8994 ( .B1(pipeline_regfile_data[1000]), .B2(n6765), .C1(
        pipeline_regfile_data[744]), .C2(n6761), .A(n8552), .ZN(n8531) );
  INV_X4 U8995 ( .A(n8553), .ZN(n8552) );
  AOI221_X2 U8996 ( .B1(pipeline_regfile_data[552]), .B2(n8299), .C1(
        pipeline_regfile_data[808]), .C2(n8300), .A(n8554), .ZN(n8553) );
  AND2_X1 U8997 ( .A1(pipeline_regfile_data[616]), .A2(n8302), .ZN(n8554) );
  NAND2_X2 U8998 ( .A1(n8556), .A2(n8557), .ZN(n8555) );
  NAND2_X2 U8999 ( .A1(pipeline_regfile_data[648]), .A2(n6769), .ZN(n8557) );
  NAND2_X2 U9000 ( .A1(pipeline_regfile_data[872]), .A2(n6770), .ZN(n8556) );
  AOI221_X2 U9001 ( .B1(pipeline_regfile_data[520]), .B2(n6709), .C1(
        pipeline_regfile_data[968]), .C2(n6763), .A(n8558), .ZN(n8529) );
  INV_X4 U9002 ( .A(n8559), .ZN(n8558) );
  AOI221_X2 U9003 ( .B1(pipeline_regfile_data[776]), .B2(n6766), .C1(
        pipeline_regfile_data[584]), .C2(n6762), .A(n8560), .ZN(n8559) );
  AND2_X1 U9004 ( .A1(pipeline_regfile_data[840]), .A2(n6768), .ZN(n8560) );
  AOI221_X2 U9005 ( .B1(pipeline_regfile_data[937]), .B2(n6767), .C1(
        pipeline_regfile_data[681]), .C2(n6764), .A(n8565), .ZN(n8564) );
  OAI22_X2 U9006 ( .A1(n8566), .A2(n8278), .B1(n8567), .B2(n9306), .ZN(n8565)
         );
  AND2_X1 U9007 ( .A1(n8568), .A2(n8569), .ZN(n8567) );
  AOI221_X2 U9008 ( .B1(pipeline_regfile_data[361]), .B2(n9309), .C1(
        pipeline_regfile_data[297]), .C2(n9315), .A(n8570), .ZN(n8569) );
  NAND2_X2 U9009 ( .A1(n8571), .A2(n8572), .ZN(n8570) );
  NAND2_X2 U9010 ( .A1(pipeline_regfile_data[489]), .A2(n9318), .ZN(n8572) );
  NAND2_X2 U9011 ( .A1(pipeline_regfile_data[425]), .A2(n9321), .ZN(n8571) );
  NAND2_X2 U9012 ( .A1(n8574), .A2(n8575), .ZN(n8573) );
  NAND2_X2 U9013 ( .A1(pipeline_regfile_data[457]), .A2(n9328), .ZN(n8575) );
  NAND2_X2 U9014 ( .A1(pipeline_regfile_data[393]), .A2(n9329), .ZN(n8574) );
  AND2_X1 U9015 ( .A1(n8576), .A2(n8577), .ZN(n8566) );
  AOI221_X2 U9016 ( .B1(pipeline_regfile_data[105]), .B2(n9308), .C1(
        pipeline_regfile_data[41]), .C2(n9315), .A(n8578), .ZN(n8577) );
  NAND2_X2 U9017 ( .A1(n8579), .A2(n8580), .ZN(n8578) );
  NAND2_X2 U9018 ( .A1(pipeline_regfile_data[233]), .A2(n9318), .ZN(n8580) );
  NAND2_X2 U9019 ( .A1(pipeline_regfile_data[169]), .A2(n9321), .ZN(n8579) );
  AOI221_X2 U9020 ( .B1(pipeline_regfile_data[73]), .B2(n9324), .C1(
        pipeline_regfile_data[9]), .C2(n9327), .A(n8581), .ZN(n8576) );
  NAND2_X2 U9021 ( .A1(n8582), .A2(n8583), .ZN(n8581) );
  NAND2_X2 U9022 ( .A1(pipeline_regfile_data[201]), .A2(n9328), .ZN(n8583) );
  NAND2_X2 U9023 ( .A1(pipeline_regfile_data[137]), .A2(n9329), .ZN(n8582) );
  AOI221_X2 U9024 ( .B1(pipeline_regfile_data[1001]), .B2(n6765), .C1(
        pipeline_regfile_data[745]), .C2(n6761), .A(n8584), .ZN(n8563) );
  INV_X4 U9025 ( .A(n8585), .ZN(n8584) );
  AOI221_X2 U9026 ( .B1(pipeline_regfile_data[553]), .B2(n8299), .C1(
        pipeline_regfile_data[809]), .C2(n8300), .A(n8586), .ZN(n8585) );
  AND2_X1 U9027 ( .A1(pipeline_regfile_data[617]), .A2(n8302), .ZN(n8586) );
  NAND2_X2 U9028 ( .A1(n8588), .A2(n8589), .ZN(n8587) );
  NAND2_X2 U9029 ( .A1(pipeline_regfile_data[649]), .A2(n6769), .ZN(n8589) );
  NAND2_X2 U9030 ( .A1(pipeline_regfile_data[873]), .A2(n6770), .ZN(n8588) );
  AOI221_X2 U9031 ( .B1(pipeline_regfile_data[521]), .B2(n6709), .C1(
        pipeline_regfile_data[969]), .C2(n6763), .A(n8590), .ZN(n8561) );
  INV_X4 U9032 ( .A(n8591), .ZN(n8590) );
  AOI221_X2 U9033 ( .B1(pipeline_regfile_data[777]), .B2(n6766), .C1(
        pipeline_regfile_data[585]), .C2(n6762), .A(n8592), .ZN(n8591) );
  AND2_X1 U9034 ( .A1(pipeline_regfile_data[841]), .A2(n6768), .ZN(n8592) );
  AOI221_X2 U9035 ( .B1(pipeline_regfile_data[938]), .B2(n6767), .C1(
        pipeline_regfile_data[682]), .C2(n6764), .A(n8597), .ZN(n8596) );
  OAI22_X2 U9036 ( .A1(n8598), .A2(n8278), .B1(n8599), .B2(n9306), .ZN(n8597)
         );
  AND2_X1 U9037 ( .A1(n8600), .A2(n8601), .ZN(n8599) );
  AOI221_X2 U9038 ( .B1(pipeline_regfile_data[362]), .B2(n9308), .C1(
        pipeline_regfile_data[298]), .C2(n9315), .A(n8602), .ZN(n8601) );
  NAND2_X2 U9039 ( .A1(n8603), .A2(n8604), .ZN(n8602) );
  NAND2_X2 U9040 ( .A1(pipeline_regfile_data[490]), .A2(n9318), .ZN(n8604) );
  NAND2_X2 U9041 ( .A1(pipeline_regfile_data[426]), .A2(n9321), .ZN(n8603) );
  NAND2_X2 U9042 ( .A1(n8606), .A2(n8607), .ZN(n8605) );
  NAND2_X2 U9043 ( .A1(pipeline_regfile_data[458]), .A2(n9328), .ZN(n8607) );
  NAND2_X2 U9044 ( .A1(pipeline_regfile_data[394]), .A2(n9330), .ZN(n8606) );
  AND2_X1 U9045 ( .A1(n8608), .A2(n8609), .ZN(n8598) );
  AOI221_X2 U9046 ( .B1(pipeline_regfile_data[106]), .B2(n9309), .C1(
        pipeline_regfile_data[42]), .C2(n9315), .A(n8610), .ZN(n8609) );
  NAND2_X2 U9047 ( .A1(n8611), .A2(n8612), .ZN(n8610) );
  NAND2_X2 U9048 ( .A1(pipeline_regfile_data[234]), .A2(n9318), .ZN(n8612) );
  NAND2_X2 U9049 ( .A1(pipeline_regfile_data[170]), .A2(n9321), .ZN(n8611) );
  AOI221_X2 U9050 ( .B1(pipeline_regfile_data[74]), .B2(n9324), .C1(
        pipeline_regfile_data[10]), .C2(n9327), .A(n8613), .ZN(n8608) );
  NAND2_X2 U9051 ( .A1(n8614), .A2(n8615), .ZN(n8613) );
  NAND2_X2 U9052 ( .A1(pipeline_regfile_data[202]), .A2(n9328), .ZN(n8615) );
  NAND2_X2 U9053 ( .A1(pipeline_regfile_data[138]), .A2(n9329), .ZN(n8614) );
  AOI221_X2 U9054 ( .B1(pipeline_regfile_data[1002]), .B2(n6765), .C1(
        pipeline_regfile_data[746]), .C2(n6761), .A(n8616), .ZN(n8595) );
  INV_X4 U9055 ( .A(n8617), .ZN(n8616) );
  AOI221_X2 U9056 ( .B1(pipeline_regfile_data[554]), .B2(n8299), .C1(
        pipeline_regfile_data[810]), .C2(n8300), .A(n8618), .ZN(n8617) );
  AND2_X1 U9057 ( .A1(pipeline_regfile_data[618]), .A2(n8302), .ZN(n8618) );
  NAND2_X2 U9058 ( .A1(n8620), .A2(n8621), .ZN(n8619) );
  NAND2_X2 U9059 ( .A1(pipeline_regfile_data[650]), .A2(n6769), .ZN(n8621) );
  NAND2_X2 U9060 ( .A1(pipeline_regfile_data[874]), .A2(n6770), .ZN(n8620) );
  AOI221_X2 U9061 ( .B1(pipeline_regfile_data[522]), .B2(n6709), .C1(
        pipeline_regfile_data[970]), .C2(n6763), .A(n8622), .ZN(n8593) );
  INV_X4 U9062 ( .A(n8623), .ZN(n8622) );
  AOI221_X2 U9063 ( .B1(pipeline_regfile_data[778]), .B2(n6766), .C1(
        pipeline_regfile_data[586]), .C2(n6762), .A(n8624), .ZN(n8623) );
  AND2_X1 U9064 ( .A1(pipeline_regfile_data[842]), .A2(n6768), .ZN(n8624) );
  AOI221_X2 U9065 ( .B1(pipeline_regfile_data[939]), .B2(n6767), .C1(
        pipeline_regfile_data[683]), .C2(n6764), .A(n8629), .ZN(n8628) );
  OAI22_X2 U9066 ( .A1(n8630), .A2(n8278), .B1(n8631), .B2(n9306), .ZN(n8629)
         );
  AOI221_X2 U9067 ( .B1(pipeline_regfile_data[363]), .B2(n9309), .C1(
        pipeline_regfile_data[299]), .C2(n9315), .A(n8634), .ZN(n8633) );
  NAND2_X2 U9068 ( .A1(n8635), .A2(n8636), .ZN(n8634) );
  NAND2_X2 U9069 ( .A1(pipeline_regfile_data[491]), .A2(n9318), .ZN(n8636) );
  NAND2_X2 U9070 ( .A1(pipeline_regfile_data[427]), .A2(n9321), .ZN(n8635) );
  AOI221_X2 U9071 ( .B1(pipeline_regfile_data[331]), .B2(n9324), .C1(
        pipeline_regfile_data[267]), .C2(n9327), .A(n8637), .ZN(n8632) );
  NAND2_X2 U9072 ( .A1(n8638), .A2(n8639), .ZN(n8637) );
  NAND2_X2 U9073 ( .A1(pipeline_regfile_data[459]), .A2(n9328), .ZN(n8639) );
  NAND2_X2 U9074 ( .A1(pipeline_regfile_data[395]), .A2(n9329), .ZN(n8638) );
  AND2_X1 U9075 ( .A1(n8640), .A2(n8641), .ZN(n8630) );
  AOI221_X2 U9076 ( .B1(pipeline_regfile_data[107]), .B2(n9308), .C1(
        pipeline_regfile_data[43]), .C2(n9315), .A(n8642), .ZN(n8641) );
  NAND2_X2 U9077 ( .A1(n8643), .A2(n8644), .ZN(n8642) );
  NAND2_X2 U9078 ( .A1(pipeline_regfile_data[235]), .A2(n9318), .ZN(n8644) );
  NAND2_X2 U9079 ( .A1(pipeline_regfile_data[171]), .A2(n9321), .ZN(n8643) );
  AOI221_X2 U9080 ( .B1(pipeline_regfile_data[75]), .B2(n9324), .C1(
        pipeline_regfile_data[11]), .C2(n9327), .A(n8645), .ZN(n8640) );
  NAND2_X2 U9081 ( .A1(n8646), .A2(n8647), .ZN(n8645) );
  NAND2_X2 U9082 ( .A1(pipeline_regfile_data[203]), .A2(n9328), .ZN(n8647) );
  NAND2_X2 U9083 ( .A1(pipeline_regfile_data[139]), .A2(n9329), .ZN(n8646) );
  AOI221_X2 U9084 ( .B1(pipeline_regfile_data[1003]), .B2(n6765), .C1(
        pipeline_regfile_data[747]), .C2(n6761), .A(n8648), .ZN(n8627) );
  INV_X4 U9085 ( .A(n8649), .ZN(n8648) );
  AOI221_X2 U9086 ( .B1(pipeline_regfile_data[555]), .B2(n8299), .C1(
        pipeline_regfile_data[811]), .C2(n8300), .A(n8650), .ZN(n8649) );
  AND2_X1 U9087 ( .A1(pipeline_regfile_data[619]), .A2(n8302), .ZN(n8650) );
  NAND2_X2 U9088 ( .A1(n8652), .A2(n8653), .ZN(n8651) );
  NAND2_X2 U9089 ( .A1(pipeline_regfile_data[651]), .A2(n6769), .ZN(n8653) );
  NAND2_X2 U9090 ( .A1(pipeline_regfile_data[875]), .A2(n6770), .ZN(n8652) );
  AOI221_X2 U9091 ( .B1(pipeline_regfile_data[523]), .B2(n6709), .C1(
        pipeline_regfile_data[971]), .C2(n6763), .A(n8654), .ZN(n8625) );
  INV_X4 U9092 ( .A(n8655), .ZN(n8654) );
  AOI221_X2 U9093 ( .B1(pipeline_regfile_data[779]), .B2(n6766), .C1(
        pipeline_regfile_data[587]), .C2(n6762), .A(n8656), .ZN(n8655) );
  AND2_X1 U9094 ( .A1(pipeline_regfile_data[843]), .A2(n6768), .ZN(n8656) );
  AOI221_X2 U9095 ( .B1(pipeline_regfile_data[940]), .B2(n6767), .C1(
        pipeline_regfile_data[684]), .C2(n6764), .A(n8661), .ZN(n8660) );
  OAI22_X2 U9096 ( .A1(n8662), .A2(n8278), .B1(n8663), .B2(n9306), .ZN(n8661)
         );
  AND2_X1 U9097 ( .A1(n8664), .A2(n8665), .ZN(n8663) );
  AOI221_X2 U9098 ( .B1(pipeline_regfile_data[364]), .B2(n9308), .C1(
        pipeline_regfile_data[300]), .C2(n9315), .A(n8666), .ZN(n8665) );
  NAND2_X2 U9099 ( .A1(n8667), .A2(n8668), .ZN(n8666) );
  NAND2_X2 U9100 ( .A1(pipeline_regfile_data[492]), .A2(n9318), .ZN(n8668) );
  NAND2_X2 U9101 ( .A1(pipeline_regfile_data[428]), .A2(n9321), .ZN(n8667) );
  AOI221_X2 U9102 ( .B1(pipeline_regfile_data[332]), .B2(n9324), .C1(
        pipeline_regfile_data[268]), .C2(n9327), .A(n8669), .ZN(n8664) );
  NAND2_X2 U9103 ( .A1(n8670), .A2(n8671), .ZN(n8669) );
  NAND2_X2 U9104 ( .A1(pipeline_regfile_data[460]), .A2(n9328), .ZN(n8671) );
  NAND2_X2 U9105 ( .A1(pipeline_regfile_data[396]), .A2(n9330), .ZN(n8670) );
  AND2_X1 U9106 ( .A1(n8672), .A2(n8673), .ZN(n8662) );
  AOI221_X2 U9107 ( .B1(pipeline_regfile_data[108]), .B2(n9308), .C1(
        pipeline_regfile_data[44]), .C2(n9315), .A(n8674), .ZN(n8673) );
  NAND2_X2 U9108 ( .A1(n8675), .A2(n8676), .ZN(n8674) );
  NAND2_X2 U9109 ( .A1(pipeline_regfile_data[236]), .A2(n9318), .ZN(n8676) );
  NAND2_X2 U9110 ( .A1(pipeline_regfile_data[172]), .A2(n9321), .ZN(n8675) );
  AOI221_X2 U9111 ( .B1(pipeline_regfile_data[76]), .B2(n9324), .C1(
        pipeline_regfile_data[12]), .C2(n9327), .A(n8677), .ZN(n8672) );
  NAND2_X2 U9112 ( .A1(n8678), .A2(n8679), .ZN(n8677) );
  NAND2_X2 U9113 ( .A1(pipeline_regfile_data[204]), .A2(n9328), .ZN(n8679) );
  NAND2_X2 U9114 ( .A1(pipeline_regfile_data[140]), .A2(n9329), .ZN(n8678) );
  AOI221_X2 U9115 ( .B1(pipeline_regfile_data[1004]), .B2(n6765), .C1(
        pipeline_regfile_data[748]), .C2(n6761), .A(n8680), .ZN(n8659) );
  INV_X4 U9116 ( .A(n8681), .ZN(n8680) );
  AOI221_X2 U9117 ( .B1(pipeline_regfile_data[556]), .B2(n8299), .C1(
        pipeline_regfile_data[812]), .C2(n8300), .A(n8682), .ZN(n8681) );
  AND2_X1 U9118 ( .A1(pipeline_regfile_data[620]), .A2(n8302), .ZN(n8682) );
  NAND2_X2 U9119 ( .A1(n8684), .A2(n8685), .ZN(n8683) );
  NAND2_X2 U9120 ( .A1(pipeline_regfile_data[652]), .A2(n6769), .ZN(n8685) );
  NAND2_X2 U9121 ( .A1(pipeline_regfile_data[876]), .A2(n6770), .ZN(n8684) );
  AOI221_X2 U9122 ( .B1(pipeline_regfile_data[524]), .B2(n6709), .C1(
        pipeline_regfile_data[972]), .C2(n6763), .A(n8686), .ZN(n8657) );
  INV_X4 U9123 ( .A(n8687), .ZN(n8686) );
  AOI221_X2 U9124 ( .B1(pipeline_regfile_data[780]), .B2(n6766), .C1(
        pipeline_regfile_data[588]), .C2(n6762), .A(n8688), .ZN(n8687) );
  AND2_X1 U9125 ( .A1(pipeline_regfile_data[844]), .A2(n6768), .ZN(n8688) );
  AOI221_X2 U9126 ( .B1(pipeline_regfile_data[941]), .B2(n6767), .C1(
        pipeline_regfile_data[685]), .C2(n6764), .A(n8693), .ZN(n8692) );
  OAI22_X2 U9127 ( .A1(n8694), .A2(n8278), .B1(n8695), .B2(n9306), .ZN(n8693)
         );
  NAND2_X2 U9128 ( .A1(n8699), .A2(n8700), .ZN(n8698) );
  NAND2_X2 U9129 ( .A1(pipeline_regfile_data[493]), .A2(n9318), .ZN(n8700) );
  NAND2_X2 U9130 ( .A1(pipeline_regfile_data[429]), .A2(n9321), .ZN(n8699) );
  AOI221_X2 U9131 ( .B1(pipeline_regfile_data[333]), .B2(n9324), .C1(
        pipeline_regfile_data[269]), .C2(n9326), .A(n8701), .ZN(n8696) );
  NAND2_X2 U9132 ( .A1(n8702), .A2(n8703), .ZN(n8701) );
  NAND2_X2 U9133 ( .A1(pipeline_regfile_data[461]), .A2(n9328), .ZN(n8703) );
  NAND2_X2 U9134 ( .A1(pipeline_regfile_data[397]), .A2(n9330), .ZN(n8702) );
  AND2_X1 U9135 ( .A1(n8704), .A2(n8705), .ZN(n8694) );
  NAND2_X2 U9136 ( .A1(n8707), .A2(n8708), .ZN(n8706) );
  NAND2_X2 U9137 ( .A1(pipeline_regfile_data[237]), .A2(n9319), .ZN(n8708) );
  NAND2_X2 U9138 ( .A1(pipeline_regfile_data[173]), .A2(n9321), .ZN(n8707) );
  AOI221_X2 U9139 ( .B1(pipeline_regfile_data[77]), .B2(n9324), .C1(
        pipeline_regfile_data[13]), .C2(n9326), .A(n8709), .ZN(n8704) );
  NAND2_X2 U9140 ( .A1(n8710), .A2(n8711), .ZN(n8709) );
  NAND2_X2 U9141 ( .A1(pipeline_regfile_data[205]), .A2(n9328), .ZN(n8711) );
  NAND2_X2 U9142 ( .A1(pipeline_regfile_data[141]), .A2(n9329), .ZN(n8710) );
  AOI221_X2 U9143 ( .B1(pipeline_regfile_data[1005]), .B2(n6765), .C1(
        pipeline_regfile_data[749]), .C2(n6761), .A(n8712), .ZN(n8691) );
  INV_X4 U9144 ( .A(n8713), .ZN(n8712) );
  AOI221_X2 U9145 ( .B1(pipeline_regfile_data[557]), .B2(n8299), .C1(
        pipeline_regfile_data[813]), .C2(n8300), .A(n8714), .ZN(n8713) );
  AND2_X1 U9146 ( .A1(pipeline_regfile_data[621]), .A2(n8302), .ZN(n8714) );
  AOI221_X2 U9147 ( .B1(pipeline_regfile_data[717]), .B2(n6773), .C1(
        pipeline_regfile_data[909]), .C2(n6772), .A(n8715), .ZN(n8690) );
  NAND2_X2 U9148 ( .A1(n8716), .A2(n8717), .ZN(n8715) );
  NAND2_X2 U9149 ( .A1(pipeline_regfile_data[653]), .A2(n6769), .ZN(n8717) );
  NAND2_X2 U9150 ( .A1(pipeline_regfile_data[877]), .A2(n6770), .ZN(n8716) );
  INV_X4 U9151 ( .A(n8719), .ZN(n8718) );
  AOI221_X2 U9152 ( .B1(pipeline_regfile_data[781]), .B2(n6766), .C1(
        pipeline_regfile_data[589]), .C2(n6762), .A(n8720), .ZN(n8719) );
  AND2_X1 U9153 ( .A1(pipeline_regfile_data[845]), .A2(n6768), .ZN(n8720) );
  AOI221_X2 U9154 ( .B1(pipeline_regfile_data[942]), .B2(n6767), .C1(
        pipeline_regfile_data[686]), .C2(n6764), .A(n8725), .ZN(n8724) );
  OAI22_X2 U9155 ( .A1(n8726), .A2(n8278), .B1(n8727), .B2(n9306), .ZN(n8725)
         );
  AND2_X1 U9156 ( .A1(n8728), .A2(n8729), .ZN(n8727) );
  AOI221_X2 U9157 ( .B1(pipeline_regfile_data[366]), .B2(n9309), .C1(
        pipeline_regfile_data[302]), .C2(n9314), .A(n8730), .ZN(n8729) );
  NAND2_X2 U9158 ( .A1(n8731), .A2(n8732), .ZN(n8730) );
  NAND2_X2 U9159 ( .A1(pipeline_regfile_data[494]), .A2(n9319), .ZN(n8732) );
  NAND2_X2 U9160 ( .A1(pipeline_regfile_data[430]), .A2(n9321), .ZN(n8731) );
  AOI221_X2 U9161 ( .B1(pipeline_regfile_data[334]), .B2(n9325), .C1(
        pipeline_regfile_data[270]), .C2(n9326), .A(n8733), .ZN(n8728) );
  NAND2_X2 U9162 ( .A1(n8734), .A2(n8735), .ZN(n8733) );
  NAND2_X2 U9163 ( .A1(pipeline_regfile_data[462]), .A2(n9328), .ZN(n8735) );
  NAND2_X2 U9164 ( .A1(pipeline_regfile_data[398]), .A2(n9329), .ZN(n8734) );
  AND2_X1 U9165 ( .A1(n8736), .A2(n8737), .ZN(n8726) );
  AOI221_X2 U9166 ( .B1(pipeline_regfile_data[110]), .B2(n9309), .C1(
        pipeline_regfile_data[46]), .C2(n9313), .A(n8738), .ZN(n8737) );
  NAND2_X2 U9167 ( .A1(n8739), .A2(n8740), .ZN(n8738) );
  NAND2_X2 U9168 ( .A1(pipeline_regfile_data[238]), .A2(n9319), .ZN(n8740) );
  NAND2_X2 U9169 ( .A1(pipeline_regfile_data[174]), .A2(n9321), .ZN(n8739) );
  AOI221_X2 U9170 ( .B1(pipeline_regfile_data[78]), .B2(n9324), .C1(
        pipeline_regfile_data[14]), .C2(n9326), .A(n8741), .ZN(n8736) );
  NAND2_X2 U9171 ( .A1(n8742), .A2(n8743), .ZN(n8741) );
  NAND2_X2 U9172 ( .A1(pipeline_regfile_data[206]), .A2(n9328), .ZN(n8743) );
  NAND2_X2 U9173 ( .A1(pipeline_regfile_data[142]), .A2(n9332), .ZN(n8742) );
  AOI221_X2 U9174 ( .B1(pipeline_regfile_data[1006]), .B2(n6765), .C1(
        pipeline_regfile_data[750]), .C2(n6761), .A(n8744), .ZN(n8723) );
  INV_X4 U9175 ( .A(n8745), .ZN(n8744) );
  AOI221_X2 U9176 ( .B1(pipeline_regfile_data[558]), .B2(n8299), .C1(
        pipeline_regfile_data[814]), .C2(n8300), .A(n8746), .ZN(n8745) );
  AND2_X1 U9177 ( .A1(pipeline_regfile_data[622]), .A2(n8302), .ZN(n8746) );
  NAND2_X2 U9178 ( .A1(n8748), .A2(n8749), .ZN(n8747) );
  NAND2_X2 U9179 ( .A1(pipeline_regfile_data[654]), .A2(n6769), .ZN(n8749) );
  NAND2_X2 U9180 ( .A1(pipeline_regfile_data[878]), .A2(n6770), .ZN(n8748) );
  AOI221_X2 U9181 ( .B1(pipeline_regfile_data[526]), .B2(n6709), .C1(
        pipeline_regfile_data[974]), .C2(n6763), .A(n8750), .ZN(n8721) );
  INV_X4 U9182 ( .A(n8751), .ZN(n8750) );
  AOI221_X2 U9183 ( .B1(pipeline_regfile_data[782]), .B2(n6766), .C1(
        pipeline_regfile_data[590]), .C2(n6762), .A(n8752), .ZN(n8751) );
  AND2_X1 U9184 ( .A1(pipeline_regfile_data[846]), .A2(n6768), .ZN(n8752) );
  AOI221_X2 U9185 ( .B1(pipeline_regfile_data[943]), .B2(n6767), .C1(
        pipeline_regfile_data[687]), .C2(n6764), .A(n8757), .ZN(n8756) );
  OAI22_X2 U9186 ( .A1(n8758), .A2(n8278), .B1(n8759), .B2(n9306), .ZN(n8757)
         );
  AND2_X1 U9187 ( .A1(n8760), .A2(n8761), .ZN(n8759) );
  NAND2_X2 U9188 ( .A1(n8763), .A2(n8764), .ZN(n8762) );
  NAND2_X2 U9189 ( .A1(pipeline_regfile_data[495]), .A2(n9319), .ZN(n8764) );
  NAND2_X2 U9190 ( .A1(pipeline_regfile_data[431]), .A2(n9321), .ZN(n8763) );
  AOI221_X2 U9191 ( .B1(pipeline_regfile_data[335]), .B2(n9324), .C1(
        pipeline_regfile_data[271]), .C2(n9326), .A(n8765), .ZN(n8760) );
  NAND2_X2 U9192 ( .A1(n8766), .A2(n8767), .ZN(n8765) );
  NAND2_X2 U9193 ( .A1(pipeline_regfile_data[463]), .A2(n9328), .ZN(n8767) );
  NAND2_X2 U9194 ( .A1(pipeline_regfile_data[399]), .A2(n9329), .ZN(n8766) );
  AND2_X1 U9195 ( .A1(n8768), .A2(n8769), .ZN(n8758) );
  AOI221_X2 U9196 ( .B1(pipeline_regfile_data[111]), .B2(n9309), .C1(
        pipeline_regfile_data[47]), .C2(n9314), .A(n8770), .ZN(n8769) );
  NAND2_X2 U9197 ( .A1(n8771), .A2(n8772), .ZN(n8770) );
  NAND2_X2 U9198 ( .A1(pipeline_regfile_data[239]), .A2(n9319), .ZN(n8772) );
  NAND2_X2 U9199 ( .A1(pipeline_regfile_data[175]), .A2(n9321), .ZN(n8771) );
  AOI221_X2 U9200 ( .B1(pipeline_regfile_data[79]), .B2(n9325), .C1(
        pipeline_regfile_data[15]), .C2(n9326), .A(n8773), .ZN(n8768) );
  NAND2_X2 U9201 ( .A1(n8774), .A2(n8775), .ZN(n8773) );
  NAND2_X2 U9202 ( .A1(pipeline_regfile_data[207]), .A2(n9328), .ZN(n8775) );
  NAND2_X2 U9203 ( .A1(pipeline_regfile_data[143]), .A2(n9332), .ZN(n8774) );
  AOI221_X2 U9204 ( .B1(pipeline_regfile_data[1007]), .B2(n6765), .C1(
        pipeline_regfile_data[751]), .C2(n6761), .A(n8776), .ZN(n8755) );
  INV_X4 U9205 ( .A(n8777), .ZN(n8776) );
  AOI221_X2 U9206 ( .B1(pipeline_regfile_data[559]), .B2(n8299), .C1(
        pipeline_regfile_data[815]), .C2(n8300), .A(n8778), .ZN(n8777) );
  AND2_X1 U9207 ( .A1(pipeline_regfile_data[623]), .A2(n8302), .ZN(n8778) );
  NAND2_X2 U9208 ( .A1(n8780), .A2(n8781), .ZN(n8779) );
  NAND2_X2 U9209 ( .A1(pipeline_regfile_data[655]), .A2(n6769), .ZN(n8781) );
  NAND2_X2 U9210 ( .A1(pipeline_regfile_data[879]), .A2(n6770), .ZN(n8780) );
  AOI221_X2 U9211 ( .B1(pipeline_regfile_data[527]), .B2(n6709), .C1(
        pipeline_regfile_data[975]), .C2(n6763), .A(n8782), .ZN(n8753) );
  INV_X4 U9212 ( .A(n8783), .ZN(n8782) );
  AOI221_X2 U9213 ( .B1(pipeline_regfile_data[783]), .B2(n6766), .C1(
        pipeline_regfile_data[591]), .C2(n6762), .A(n8784), .ZN(n8783) );
  AND2_X1 U9214 ( .A1(pipeline_regfile_data[847]), .A2(n6768), .ZN(n8784) );
  AOI221_X2 U9215 ( .B1(pipeline_regfile_data[944]), .B2(n6767), .C1(
        pipeline_regfile_data[688]), .C2(n6764), .A(n8789), .ZN(n8788) );
  OAI22_X2 U9216 ( .A1(n8790), .A2(n8278), .B1(n8791), .B2(n9306), .ZN(n8789)
         );
  NAND2_X2 U9217 ( .A1(n8795), .A2(n8796), .ZN(n8794) );
  NAND2_X2 U9218 ( .A1(pipeline_regfile_data[496]), .A2(n9319), .ZN(n8796) );
  NAND2_X2 U9219 ( .A1(pipeline_regfile_data[432]), .A2(n9321), .ZN(n8795) );
  AOI221_X2 U9220 ( .B1(pipeline_regfile_data[336]), .B2(n9325), .C1(
        pipeline_regfile_data[272]), .C2(n9326), .A(n8797), .ZN(n8792) );
  NAND2_X2 U9221 ( .A1(n8798), .A2(n8799), .ZN(n8797) );
  NAND2_X2 U9222 ( .A1(pipeline_regfile_data[464]), .A2(n9328), .ZN(n8799) );
  NAND2_X2 U9223 ( .A1(pipeline_regfile_data[400]), .A2(n9331), .ZN(n8798) );
  AND2_X1 U9224 ( .A1(n8800), .A2(n8801), .ZN(n8790) );
  NAND2_X2 U9225 ( .A1(n8803), .A2(n8804), .ZN(n8802) );
  NAND2_X2 U9226 ( .A1(pipeline_regfile_data[240]), .A2(n9319), .ZN(n8804) );
  NAND2_X2 U9227 ( .A1(pipeline_regfile_data[176]), .A2(n9321), .ZN(n8803) );
  AOI221_X2 U9228 ( .B1(pipeline_regfile_data[80]), .B2(n9325), .C1(
        pipeline_regfile_data[16]), .C2(n9326), .A(n8805), .ZN(n8800) );
  NAND2_X2 U9229 ( .A1(n8806), .A2(n8807), .ZN(n8805) );
  NAND2_X2 U9230 ( .A1(pipeline_regfile_data[208]), .A2(n9328), .ZN(n8807) );
  NAND2_X2 U9231 ( .A1(pipeline_regfile_data[144]), .A2(n9331), .ZN(n8806) );
  AOI221_X2 U9232 ( .B1(pipeline_regfile_data[1008]), .B2(n6765), .C1(
        pipeline_regfile_data[752]), .C2(n6761), .A(n8808), .ZN(n8787) );
  INV_X4 U9233 ( .A(n8809), .ZN(n8808) );
  AOI221_X2 U9234 ( .B1(pipeline_regfile_data[560]), .B2(n8299), .C1(
        pipeline_regfile_data[816]), .C2(n8300), .A(n8810), .ZN(n8809) );
  AND2_X1 U9235 ( .A1(pipeline_regfile_data[624]), .A2(n8302), .ZN(n8810) );
  AOI221_X2 U9236 ( .B1(pipeline_regfile_data[720]), .B2(n6773), .C1(
        pipeline_regfile_data[912]), .C2(n6772), .A(n8811), .ZN(n8786) );
  NAND2_X2 U9237 ( .A1(n8812), .A2(n8813), .ZN(n8811) );
  NAND2_X2 U9238 ( .A1(pipeline_regfile_data[656]), .A2(n6769), .ZN(n8813) );
  NAND2_X2 U9239 ( .A1(pipeline_regfile_data[880]), .A2(n6770), .ZN(n8812) );
  AOI221_X2 U9240 ( .B1(pipeline_regfile_data[528]), .B2(n6709), .C1(
        pipeline_regfile_data[976]), .C2(n6763), .A(n8814), .ZN(n8785) );
  INV_X4 U9241 ( .A(n8815), .ZN(n8814) );
  AOI221_X2 U9242 ( .B1(pipeline_regfile_data[784]), .B2(n6766), .C1(
        pipeline_regfile_data[592]), .C2(n6762), .A(n8816), .ZN(n8815) );
  AND2_X1 U9243 ( .A1(pipeline_regfile_data[848]), .A2(n6768), .ZN(n8816) );
  AOI221_X2 U9244 ( .B1(pipeline_regfile_data[945]), .B2(n6767), .C1(
        pipeline_regfile_data[689]), .C2(n6764), .A(n8821), .ZN(n8820) );
  OAI22_X2 U9245 ( .A1(n8822), .A2(n8278), .B1(n8823), .B2(n9306), .ZN(n8821)
         );
  AND2_X1 U9246 ( .A1(n8824), .A2(n8825), .ZN(n8823) );
  NAND2_X2 U9247 ( .A1(n8827), .A2(n8828), .ZN(n8826) );
  NAND2_X2 U9248 ( .A1(pipeline_regfile_data[497]), .A2(n9319), .ZN(n8828) );
  NAND2_X2 U9249 ( .A1(pipeline_regfile_data[433]), .A2(n9321), .ZN(n8827) );
  AOI221_X2 U9250 ( .B1(pipeline_regfile_data[337]), .B2(n9325), .C1(
        pipeline_regfile_data[273]), .C2(n9326), .A(n8829), .ZN(n8824) );
  NAND2_X2 U9251 ( .A1(n8830), .A2(n8831), .ZN(n8829) );
  NAND2_X2 U9252 ( .A1(pipeline_regfile_data[465]), .A2(n9328), .ZN(n8831) );
  NAND2_X2 U9253 ( .A1(pipeline_regfile_data[401]), .A2(n9330), .ZN(n8830) );
  AND2_X1 U9254 ( .A1(n8832), .A2(n8833), .ZN(n8822) );
  AOI221_X2 U9255 ( .B1(pipeline_regfile_data[113]), .B2(n9309), .C1(
        pipeline_regfile_data[49]), .C2(n9313), .A(n8834), .ZN(n8833) );
  NAND2_X2 U9256 ( .A1(n8835), .A2(n8836), .ZN(n8834) );
  NAND2_X2 U9257 ( .A1(pipeline_regfile_data[241]), .A2(n9319), .ZN(n8836) );
  NAND2_X2 U9258 ( .A1(pipeline_regfile_data[177]), .A2(n9321), .ZN(n8835) );
  AOI221_X2 U9259 ( .B1(pipeline_regfile_data[81]), .B2(n9325), .C1(
        pipeline_regfile_data[17]), .C2(n9326), .A(n8837), .ZN(n8832) );
  NAND2_X2 U9260 ( .A1(n8838), .A2(n8839), .ZN(n8837) );
  NAND2_X2 U9261 ( .A1(pipeline_regfile_data[209]), .A2(n9328), .ZN(n8839) );
  NAND2_X2 U9262 ( .A1(pipeline_regfile_data[145]), .A2(n9329), .ZN(n8838) );
  AOI221_X2 U9263 ( .B1(pipeline_regfile_data[1009]), .B2(n6765), .C1(
        pipeline_regfile_data[753]), .C2(n6761), .A(n8840), .ZN(n8819) );
  INV_X4 U9264 ( .A(n8841), .ZN(n8840) );
  AOI221_X2 U9265 ( .B1(pipeline_regfile_data[561]), .B2(n8299), .C1(
        pipeline_regfile_data[817]), .C2(n8300), .A(n8842), .ZN(n8841) );
  AND2_X1 U9266 ( .A1(pipeline_regfile_data[625]), .A2(n8302), .ZN(n8842) );
  NAND2_X2 U9267 ( .A1(n8844), .A2(n8845), .ZN(n8843) );
  NAND2_X2 U9268 ( .A1(pipeline_regfile_data[657]), .A2(n6769), .ZN(n8845) );
  NAND2_X2 U9269 ( .A1(pipeline_regfile_data[881]), .A2(n6770), .ZN(n8844) );
  AOI221_X2 U9270 ( .B1(pipeline_regfile_data[529]), .B2(n6709), .C1(
        pipeline_regfile_data[977]), .C2(n6763), .A(n8846), .ZN(n8817) );
  INV_X4 U9271 ( .A(n8847), .ZN(n8846) );
  AOI221_X2 U9272 ( .B1(pipeline_regfile_data[785]), .B2(n6766), .C1(
        pipeline_regfile_data[593]), .C2(n6762), .A(n8848), .ZN(n8847) );
  AND2_X1 U9273 ( .A1(pipeline_regfile_data[849]), .A2(n6768), .ZN(n8848) );
  AOI221_X2 U9274 ( .B1(pipeline_regfile_data[946]), .B2(n6767), .C1(
        pipeline_regfile_data[690]), .C2(n6764), .A(n8853), .ZN(n8852) );
  OAI22_X2 U9275 ( .A1(n8854), .A2(n8278), .B1(n8855), .B2(n9306), .ZN(n8853)
         );
  AND2_X1 U9276 ( .A1(n8856), .A2(n8857), .ZN(n8855) );
  NAND2_X2 U9277 ( .A1(n8859), .A2(n8860), .ZN(n8858) );
  NAND2_X2 U9278 ( .A1(pipeline_regfile_data[498]), .A2(n9319), .ZN(n8860) );
  NAND2_X2 U9279 ( .A1(pipeline_regfile_data[434]), .A2(n9321), .ZN(n8859) );
  AOI221_X2 U9280 ( .B1(pipeline_regfile_data[338]), .B2(n9324), .C1(
        pipeline_regfile_data[274]), .C2(n9326), .A(n8861), .ZN(n8856) );
  NAND2_X2 U9281 ( .A1(n8862), .A2(n8863), .ZN(n8861) );
  NAND2_X2 U9282 ( .A1(pipeline_regfile_data[466]), .A2(n9328), .ZN(n8863) );
  NAND2_X2 U9283 ( .A1(pipeline_regfile_data[402]), .A2(n9330), .ZN(n8862) );
  AND2_X1 U9284 ( .A1(n8864), .A2(n8865), .ZN(n8854) );
  AOI221_X2 U9285 ( .B1(pipeline_regfile_data[114]), .B2(n9309), .C1(
        pipeline_regfile_data[50]), .C2(n9313), .A(n8866), .ZN(n8865) );
  NAND2_X2 U9286 ( .A1(n8867), .A2(n8868), .ZN(n8866) );
  NAND2_X2 U9287 ( .A1(pipeline_regfile_data[242]), .A2(n9319), .ZN(n8868) );
  NAND2_X2 U9288 ( .A1(pipeline_regfile_data[178]), .A2(n9321), .ZN(n8867) );
  AOI221_X2 U9289 ( .B1(pipeline_regfile_data[82]), .B2(n9325), .C1(
        pipeline_regfile_data[18]), .C2(n9326), .A(n8869), .ZN(n8864) );
  NAND2_X2 U9290 ( .A1(n8870), .A2(n8871), .ZN(n8869) );
  NAND2_X2 U9291 ( .A1(pipeline_regfile_data[210]), .A2(n9328), .ZN(n8871) );
  NAND2_X2 U9292 ( .A1(pipeline_regfile_data[146]), .A2(n9330), .ZN(n8870) );
  AOI221_X2 U9293 ( .B1(pipeline_regfile_data[1010]), .B2(n6765), .C1(
        pipeline_regfile_data[754]), .C2(n6761), .A(n8872), .ZN(n8851) );
  INV_X4 U9294 ( .A(n8873), .ZN(n8872) );
  AOI221_X2 U9295 ( .B1(pipeline_regfile_data[562]), .B2(n8299), .C1(
        pipeline_regfile_data[818]), .C2(n8300), .A(n8874), .ZN(n8873) );
  AND2_X1 U9296 ( .A1(pipeline_regfile_data[626]), .A2(n8302), .ZN(n8874) );
  NAND2_X2 U9297 ( .A1(n8876), .A2(n8877), .ZN(n8875) );
  NAND2_X2 U9298 ( .A1(pipeline_regfile_data[658]), .A2(n6769), .ZN(n8877) );
  NAND2_X2 U9299 ( .A1(pipeline_regfile_data[882]), .A2(n6770), .ZN(n8876) );
  AOI221_X2 U9300 ( .B1(pipeline_regfile_data[530]), .B2(n6709), .C1(
        pipeline_regfile_data[978]), .C2(n6763), .A(n8878), .ZN(n8849) );
  INV_X4 U9301 ( .A(n8879), .ZN(n8878) );
  AOI221_X2 U9302 ( .B1(pipeline_regfile_data[786]), .B2(n6766), .C1(
        pipeline_regfile_data[594]), .C2(n6762), .A(n8880), .ZN(n8879) );
  AND2_X1 U9303 ( .A1(pipeline_regfile_data[850]), .A2(n6768), .ZN(n8880) );
  AOI221_X2 U9304 ( .B1(pipeline_regfile_data[947]), .B2(n6767), .C1(
        pipeline_regfile_data[691]), .C2(n6764), .A(n8885), .ZN(n8884) );
  OAI22_X2 U9305 ( .A1(n8886), .A2(n8278), .B1(n8887), .B2(n9306), .ZN(n8885)
         );
  NAND2_X2 U9306 ( .A1(n8891), .A2(n8892), .ZN(n8890) );
  NAND2_X2 U9307 ( .A1(pipeline_regfile_data[499]), .A2(n9319), .ZN(n8892) );
  NAND2_X2 U9308 ( .A1(pipeline_regfile_data[435]), .A2(n9321), .ZN(n8891) );
  AOI221_X2 U9309 ( .B1(pipeline_regfile_data[339]), .B2(n9324), .C1(
        pipeline_regfile_data[275]), .C2(n9326), .A(n8893), .ZN(n8888) );
  NAND2_X2 U9310 ( .A1(n8894), .A2(n8895), .ZN(n8893) );
  NAND2_X2 U9311 ( .A1(pipeline_regfile_data[467]), .A2(n9328), .ZN(n8895) );
  NAND2_X2 U9312 ( .A1(pipeline_regfile_data[403]), .A2(n9331), .ZN(n8894) );
  AND2_X1 U9313 ( .A1(n8896), .A2(n8897), .ZN(n8886) );
  NAND2_X2 U9314 ( .A1(n8899), .A2(n8900), .ZN(n8898) );
  NAND2_X2 U9315 ( .A1(pipeline_regfile_data[243]), .A2(n9319), .ZN(n8900) );
  NAND2_X2 U9316 ( .A1(pipeline_regfile_data[179]), .A2(n9321), .ZN(n8899) );
  AOI221_X2 U9317 ( .B1(pipeline_regfile_data[83]), .B2(n9323), .C1(
        pipeline_regfile_data[19]), .C2(n9327), .A(n8901), .ZN(n8896) );
  NAND2_X2 U9318 ( .A1(n8902), .A2(n8903), .ZN(n8901) );
  NAND2_X2 U9319 ( .A1(pipeline_regfile_data[211]), .A2(n9328), .ZN(n8903) );
  NAND2_X2 U9320 ( .A1(pipeline_regfile_data[147]), .A2(n9329), .ZN(n8902) );
  AOI221_X2 U9321 ( .B1(pipeline_regfile_data[1011]), .B2(n6765), .C1(
        pipeline_regfile_data[755]), .C2(n6761), .A(n8904), .ZN(n8883) );
  INV_X4 U9322 ( .A(n8905), .ZN(n8904) );
  AOI221_X2 U9323 ( .B1(pipeline_regfile_data[563]), .B2(n8299), .C1(
        pipeline_regfile_data[819]), .C2(n8300), .A(n8906), .ZN(n8905) );
  AND2_X1 U9324 ( .A1(pipeline_regfile_data[627]), .A2(n8302), .ZN(n8906) );
  NAND2_X2 U9325 ( .A1(n8908), .A2(n8909), .ZN(n8907) );
  NAND2_X2 U9326 ( .A1(pipeline_regfile_data[659]), .A2(n6769), .ZN(n8909) );
  NAND2_X2 U9327 ( .A1(pipeline_regfile_data[883]), .A2(n6770), .ZN(n8908) );
  AOI221_X2 U9328 ( .B1(pipeline_regfile_data[531]), .B2(n6709), .C1(
        pipeline_regfile_data[979]), .C2(n6763), .A(n8910), .ZN(n8881) );
  INV_X4 U9329 ( .A(n8911), .ZN(n8910) );
  AOI221_X2 U9330 ( .B1(pipeline_regfile_data[787]), .B2(n6766), .C1(
        pipeline_regfile_data[595]), .C2(n6762), .A(n8912), .ZN(n8911) );
  AND2_X1 U9331 ( .A1(pipeline_regfile_data[851]), .A2(n6768), .ZN(n8912) );
  AOI221_X2 U9332 ( .B1(pipeline_regfile_data[948]), .B2(n6767), .C1(
        pipeline_regfile_data[692]), .C2(n6764), .A(n8917), .ZN(n8916) );
  OAI22_X2 U9333 ( .A1(n8918), .A2(n9305), .B1(n8919), .B2(n9306), .ZN(n8917)
         );
  AND2_X1 U9334 ( .A1(n8920), .A2(n8921), .ZN(n8919) );
  AOI221_X2 U9335 ( .B1(pipeline_regfile_data[372]), .B2(n9308), .C1(
        pipeline_regfile_data[308]), .C2(n9314), .A(n8922), .ZN(n8921) );
  NAND2_X2 U9336 ( .A1(n8923), .A2(n8924), .ZN(n8922) );
  NAND2_X2 U9337 ( .A1(pipeline_regfile_data[500]), .A2(n9320), .ZN(n8924) );
  NAND2_X2 U9338 ( .A1(pipeline_regfile_data[436]), .A2(n9321), .ZN(n8923) );
  AOI221_X2 U9339 ( .B1(pipeline_regfile_data[340]), .B2(n9323), .C1(
        pipeline_regfile_data[276]), .C2(n9327), .A(n8925), .ZN(n8920) );
  NAND2_X2 U9340 ( .A1(n8926), .A2(n8927), .ZN(n8925) );
  NAND2_X2 U9341 ( .A1(pipeline_regfile_data[468]), .A2(n9328), .ZN(n8927) );
  NAND2_X2 U9342 ( .A1(pipeline_regfile_data[404]), .A2(n9330), .ZN(n8926) );
  AND2_X1 U9343 ( .A1(n8928), .A2(n8929), .ZN(n8918) );
  NAND2_X2 U9344 ( .A1(n8931), .A2(n8932), .ZN(n8930) );
  NAND2_X2 U9345 ( .A1(pipeline_regfile_data[244]), .A2(n9320), .ZN(n8932) );
  NAND2_X2 U9346 ( .A1(pipeline_regfile_data[180]), .A2(n9321), .ZN(n8931) );
  AOI221_X2 U9347 ( .B1(pipeline_regfile_data[84]), .B2(n9323), .C1(
        pipeline_regfile_data[20]), .C2(n9327), .A(n8933), .ZN(n8928) );
  NAND2_X2 U9348 ( .A1(n8934), .A2(n8935), .ZN(n8933) );
  NAND2_X2 U9349 ( .A1(pipeline_regfile_data[212]), .A2(n9328), .ZN(n8935) );
  NAND2_X2 U9350 ( .A1(pipeline_regfile_data[148]), .A2(n9330), .ZN(n8934) );
  AOI221_X2 U9351 ( .B1(pipeline_regfile_data[1012]), .B2(n6765), .C1(
        pipeline_regfile_data[756]), .C2(n6761), .A(n8936), .ZN(n8915) );
  INV_X4 U9352 ( .A(n8937), .ZN(n8936) );
  AOI221_X2 U9353 ( .B1(pipeline_regfile_data[564]), .B2(n8299), .C1(
        pipeline_regfile_data[820]), .C2(n8300), .A(n8938), .ZN(n8937) );
  AND2_X1 U9354 ( .A1(pipeline_regfile_data[628]), .A2(n8302), .ZN(n8938) );
  NAND2_X2 U9355 ( .A1(n8940), .A2(n8941), .ZN(n8939) );
  NAND2_X2 U9356 ( .A1(pipeline_regfile_data[660]), .A2(n6769), .ZN(n8941) );
  NAND2_X2 U9357 ( .A1(pipeline_regfile_data[884]), .A2(n6770), .ZN(n8940) );
  AOI221_X2 U9358 ( .B1(pipeline_regfile_data[532]), .B2(n6709), .C1(
        pipeline_regfile_data[980]), .C2(n6763), .A(n8942), .ZN(n8913) );
  INV_X4 U9359 ( .A(n8943), .ZN(n8942) );
  AOI221_X2 U9360 ( .B1(pipeline_regfile_data[788]), .B2(n6766), .C1(
        pipeline_regfile_data[596]), .C2(n6762), .A(n8944), .ZN(n8943) );
  AND2_X1 U9361 ( .A1(pipeline_regfile_data[852]), .A2(n6768), .ZN(n8944) );
  AOI221_X2 U9362 ( .B1(pipeline_regfile_data[949]), .B2(n6767), .C1(
        pipeline_regfile_data[693]), .C2(n6764), .A(n8949), .ZN(n8948) );
  OAI22_X2 U9363 ( .A1(n8950), .A2(n9305), .B1(n8951), .B2(n9306), .ZN(n8949)
         );
  NAND2_X2 U9364 ( .A1(n8955), .A2(n8956), .ZN(n8954) );
  NAND2_X2 U9365 ( .A1(pipeline_regfile_data[501]), .A2(n9320), .ZN(n8956) );
  NAND2_X2 U9366 ( .A1(pipeline_regfile_data[437]), .A2(n9321), .ZN(n8955) );
  AOI221_X2 U9367 ( .B1(pipeline_regfile_data[341]), .B2(n9323), .C1(
        pipeline_regfile_data[277]), .C2(n9327), .A(n8957), .ZN(n8952) );
  NAND2_X2 U9368 ( .A1(n8958), .A2(n8959), .ZN(n8957) );
  NAND2_X2 U9369 ( .A1(pipeline_regfile_data[469]), .A2(n9328), .ZN(n8959) );
  NAND2_X2 U9370 ( .A1(pipeline_regfile_data[405]), .A2(n9331), .ZN(n8958) );
  AND2_X1 U9371 ( .A1(n8960), .A2(n8961), .ZN(n8950) );
  NAND2_X2 U9372 ( .A1(n8963), .A2(n8964), .ZN(n8962) );
  NAND2_X2 U9373 ( .A1(pipeline_regfile_data[245]), .A2(n9320), .ZN(n8964) );
  NAND2_X2 U9374 ( .A1(pipeline_regfile_data[181]), .A2(n9321), .ZN(n8963) );
  AOI221_X2 U9375 ( .B1(pipeline_regfile_data[85]), .B2(n9323), .C1(
        pipeline_regfile_data[21]), .C2(n9327), .A(n8965), .ZN(n8960) );
  NAND2_X2 U9376 ( .A1(n8966), .A2(n8967), .ZN(n8965) );
  NAND2_X2 U9377 ( .A1(pipeline_regfile_data[213]), .A2(n9328), .ZN(n8967) );
  NAND2_X2 U9378 ( .A1(pipeline_regfile_data[149]), .A2(n9330), .ZN(n8966) );
  AOI221_X2 U9379 ( .B1(pipeline_regfile_data[1013]), .B2(n6765), .C1(
        pipeline_regfile_data[757]), .C2(n6761), .A(n8968), .ZN(n8947) );
  INV_X4 U9380 ( .A(n8969), .ZN(n8968) );
  AOI221_X2 U9381 ( .B1(pipeline_regfile_data[565]), .B2(n8299), .C1(
        pipeline_regfile_data[821]), .C2(n8300), .A(n8970), .ZN(n8969) );
  AND2_X1 U9382 ( .A1(pipeline_regfile_data[629]), .A2(n8302), .ZN(n8970) );
  NAND2_X2 U9383 ( .A1(n8972), .A2(n8973), .ZN(n8971) );
  NAND2_X2 U9384 ( .A1(pipeline_regfile_data[661]), .A2(n6769), .ZN(n8973) );
  NAND2_X2 U9385 ( .A1(pipeline_regfile_data[885]), .A2(n6770), .ZN(n8972) );
  AOI221_X2 U9386 ( .B1(pipeline_regfile_data[533]), .B2(n6709), .C1(
        pipeline_regfile_data[981]), .C2(n6763), .A(n8974), .ZN(n8945) );
  INV_X4 U9387 ( .A(n8975), .ZN(n8974) );
  AOI221_X2 U9388 ( .B1(pipeline_regfile_data[789]), .B2(n6766), .C1(
        pipeline_regfile_data[597]), .C2(n6762), .A(n8976), .ZN(n8975) );
  AND2_X1 U9389 ( .A1(pipeline_regfile_data[853]), .A2(n6768), .ZN(n8976) );
  AOI221_X2 U9390 ( .B1(pipeline_regfile_data[950]), .B2(n6767), .C1(
        pipeline_regfile_data[694]), .C2(n6764), .A(n8981), .ZN(n8980) );
  NAND2_X2 U9391 ( .A1(n8985), .A2(n8986), .ZN(n8984) );
  NAND2_X2 U9392 ( .A1(pipeline_regfile_data[502]), .A2(n9320), .ZN(n8986) );
  NAND2_X2 U9393 ( .A1(pipeline_regfile_data[438]), .A2(n9321), .ZN(n8985) );
  AOI221_X2 U9394 ( .B1(pipeline_regfile_data[342]), .B2(n9323), .C1(
        pipeline_regfile_data[278]), .C2(n9326), .A(n8987), .ZN(n8982) );
  NAND2_X2 U9395 ( .A1(n8988), .A2(n8989), .ZN(n8987) );
  NAND2_X2 U9396 ( .A1(pipeline_regfile_data[470]), .A2(n9328), .ZN(n8989) );
  NAND2_X2 U9397 ( .A1(pipeline_regfile_data[406]), .A2(n9332), .ZN(n8988) );
  NAND2_X2 U9398 ( .A1(n8993), .A2(n8994), .ZN(n8992) );
  NAND2_X2 U9399 ( .A1(pipeline_regfile_data[246]), .A2(n9320), .ZN(n8994) );
  NAND2_X2 U9400 ( .A1(pipeline_regfile_data[182]), .A2(n9321), .ZN(n8993) );
  NAND2_X2 U9401 ( .A1(n8996), .A2(n8997), .ZN(n8995) );
  NAND2_X2 U9402 ( .A1(pipeline_regfile_data[214]), .A2(n9328), .ZN(n8997) );
  NAND2_X2 U9403 ( .A1(pipeline_regfile_data[150]), .A2(n9330), .ZN(n8996) );
  AOI221_X2 U9404 ( .B1(pipeline_regfile_data[1014]), .B2(n6765), .C1(
        pipeline_regfile_data[758]), .C2(n6761), .A(n8998), .ZN(n8979) );
  INV_X4 U9405 ( .A(n8999), .ZN(n8998) );
  AOI221_X2 U9406 ( .B1(pipeline_regfile_data[566]), .B2(n8299), .C1(
        pipeline_regfile_data[822]), .C2(n8300), .A(n9000), .ZN(n8999) );
  AND2_X1 U9407 ( .A1(pipeline_regfile_data[630]), .A2(n8302), .ZN(n9000) );
  NAND2_X2 U9408 ( .A1(n9002), .A2(n9003), .ZN(n9001) );
  NAND2_X2 U9409 ( .A1(pipeline_regfile_data[662]), .A2(n6769), .ZN(n9003) );
  NAND2_X2 U9410 ( .A1(pipeline_regfile_data[886]), .A2(n6770), .ZN(n9002) );
  AOI221_X2 U9411 ( .B1(pipeline_regfile_data[534]), .B2(n6709), .C1(
        pipeline_regfile_data[982]), .C2(n6763), .A(n9004), .ZN(n8977) );
  INV_X4 U9412 ( .A(n9005), .ZN(n9004) );
  AOI221_X2 U9413 ( .B1(pipeline_regfile_data[790]), .B2(n6766), .C1(
        pipeline_regfile_data[598]), .C2(n6762), .A(n9006), .ZN(n9005) );
  AND2_X1 U9414 ( .A1(pipeline_regfile_data[854]), .A2(n6768), .ZN(n9006) );
  AOI221_X2 U9415 ( .B1(pipeline_regfile_data[951]), .B2(n6767), .C1(
        pipeline_regfile_data[695]), .C2(n6764), .A(n9011), .ZN(n9010) );
  OAI22_X2 U9416 ( .A1(n9012), .A2(n9305), .B1(n9013), .B2(n9306), .ZN(n9011)
         );
  NAND2_X2 U9417 ( .A1(n9017), .A2(n9018), .ZN(n9016) );
  NAND2_X2 U9418 ( .A1(pipeline_regfile_data[503]), .A2(n9320), .ZN(n9018) );
  NAND2_X2 U9419 ( .A1(pipeline_regfile_data[439]), .A2(n9321), .ZN(n9017) );
  AOI221_X2 U9420 ( .B1(pipeline_regfile_data[343]), .B2(n9323), .C1(
        pipeline_regfile_data[279]), .C2(n9327), .A(n9019), .ZN(n9014) );
  NAND2_X2 U9421 ( .A1(n9020), .A2(n9021), .ZN(n9019) );
  NAND2_X2 U9422 ( .A1(pipeline_regfile_data[471]), .A2(n9328), .ZN(n9021) );
  NAND2_X2 U9423 ( .A1(pipeline_regfile_data[407]), .A2(n9330), .ZN(n9020) );
  AND2_X1 U9424 ( .A1(n9022), .A2(n9023), .ZN(n9012) );
  NAND2_X2 U9425 ( .A1(n9025), .A2(n9026), .ZN(n9024) );
  NAND2_X2 U9426 ( .A1(pipeline_regfile_data[247]), .A2(n9320), .ZN(n9026) );
  NAND2_X2 U9427 ( .A1(pipeline_regfile_data[183]), .A2(n9321), .ZN(n9025) );
  NAND2_X2 U9428 ( .A1(n9028), .A2(n9029), .ZN(n9027) );
  NAND2_X2 U9429 ( .A1(pipeline_regfile_data[215]), .A2(n9328), .ZN(n9029) );
  NAND2_X2 U9430 ( .A1(pipeline_regfile_data[151]), .A2(n9330), .ZN(n9028) );
  AOI221_X2 U9431 ( .B1(pipeline_regfile_data[1015]), .B2(n6765), .C1(
        pipeline_regfile_data[759]), .C2(n6761), .A(n9030), .ZN(n9009) );
  INV_X4 U9432 ( .A(n9031), .ZN(n9030) );
  AOI221_X2 U9433 ( .B1(pipeline_regfile_data[567]), .B2(n8299), .C1(
        pipeline_regfile_data[823]), .C2(n8300), .A(n9032), .ZN(n9031) );
  AND2_X1 U9434 ( .A1(pipeline_regfile_data[631]), .A2(n8302), .ZN(n9032) );
  AOI221_X2 U9435 ( .B1(pipeline_regfile_data[727]), .B2(n6773), .C1(
        pipeline_regfile_data[919]), .C2(n6772), .A(n9033), .ZN(n9008) );
  NAND2_X2 U9436 ( .A1(n9034), .A2(n9035), .ZN(n9033) );
  NAND2_X2 U9437 ( .A1(pipeline_regfile_data[663]), .A2(n6769), .ZN(n9035) );
  NAND2_X2 U9438 ( .A1(pipeline_regfile_data[887]), .A2(n6770), .ZN(n9034) );
  INV_X4 U9439 ( .A(n9037), .ZN(n9036) );
  AOI221_X2 U9440 ( .B1(pipeline_regfile_data[791]), .B2(n6766), .C1(
        pipeline_regfile_data[599]), .C2(n6762), .A(n9038), .ZN(n9037) );
  AND2_X1 U9441 ( .A1(pipeline_regfile_data[855]), .A2(n6768), .ZN(n9038) );
  AOI221_X2 U9442 ( .B1(pipeline_regfile_data[952]), .B2(n6767), .C1(
        pipeline_regfile_data[696]), .C2(n6764), .A(n9043), .ZN(n9042) );
  OAI22_X2 U9443 ( .A1(n9044), .A2(n9305), .B1(n9045), .B2(n9306), .ZN(n9043)
         );
  AND2_X1 U9444 ( .A1(n9046), .A2(n9047), .ZN(n9045) );
  NAND2_X2 U9445 ( .A1(n9049), .A2(n9050), .ZN(n9048) );
  NAND2_X2 U9446 ( .A1(pipeline_regfile_data[504]), .A2(n9320), .ZN(n9050) );
  NAND2_X2 U9447 ( .A1(pipeline_regfile_data[440]), .A2(n9321), .ZN(n9049) );
  AOI221_X2 U9448 ( .B1(pipeline_regfile_data[344]), .B2(n9323), .C1(
        pipeline_regfile_data[280]), .C2(n9327), .A(n9051), .ZN(n9046) );
  NAND2_X2 U9449 ( .A1(n9052), .A2(n9053), .ZN(n9051) );
  NAND2_X2 U9450 ( .A1(pipeline_regfile_data[472]), .A2(n9328), .ZN(n9053) );
  NAND2_X2 U9451 ( .A1(pipeline_regfile_data[408]), .A2(n9331), .ZN(n9052) );
  AND2_X1 U9452 ( .A1(n9054), .A2(n9055), .ZN(n9044) );
  NAND2_X2 U9453 ( .A1(n9057), .A2(n9058), .ZN(n9056) );
  NAND2_X2 U9454 ( .A1(pipeline_regfile_data[248]), .A2(n9320), .ZN(n9058) );
  NAND2_X2 U9455 ( .A1(pipeline_regfile_data[184]), .A2(n9321), .ZN(n9057) );
  AOI221_X2 U9456 ( .B1(pipeline_regfile_data[88]), .B2(n9323), .C1(
        pipeline_regfile_data[24]), .C2(n9327), .A(n9059), .ZN(n9054) );
  NAND2_X2 U9457 ( .A1(n9060), .A2(n9061), .ZN(n9059) );
  NAND2_X2 U9458 ( .A1(pipeline_regfile_data[216]), .A2(n9328), .ZN(n9061) );
  NAND2_X2 U9459 ( .A1(pipeline_regfile_data[152]), .A2(n9330), .ZN(n9060) );
  AOI221_X2 U9460 ( .B1(pipeline_regfile_data[1016]), .B2(n6765), .C1(
        pipeline_regfile_data[760]), .C2(n6761), .A(n9062), .ZN(n9041) );
  INV_X4 U9461 ( .A(n9063), .ZN(n9062) );
  AOI221_X2 U9462 ( .B1(pipeline_regfile_data[568]), .B2(n8299), .C1(
        pipeline_regfile_data[824]), .C2(n8300), .A(n9064), .ZN(n9063) );
  AND2_X1 U9463 ( .A1(pipeline_regfile_data[632]), .A2(n8302), .ZN(n9064) );
  NAND2_X2 U9464 ( .A1(n9066), .A2(n9067), .ZN(n9065) );
  NAND2_X2 U9465 ( .A1(pipeline_regfile_data[664]), .A2(n6769), .ZN(n9067) );
  NAND2_X2 U9466 ( .A1(pipeline_regfile_data[888]), .A2(n6770), .ZN(n9066) );
  AOI221_X2 U9467 ( .B1(pipeline_regfile_data[536]), .B2(n6709), .C1(
        pipeline_regfile_data[984]), .C2(n6763), .A(n9068), .ZN(n9039) );
  INV_X4 U9468 ( .A(n9069), .ZN(n9068) );
  AOI221_X2 U9469 ( .B1(pipeline_regfile_data[792]), .B2(n6766), .C1(
        pipeline_regfile_data[600]), .C2(n6762), .A(n9070), .ZN(n9069) );
  AND2_X1 U9470 ( .A1(pipeline_regfile_data[856]), .A2(n6768), .ZN(n9070) );
  AOI221_X2 U9471 ( .B1(pipeline_regfile_data[953]), .B2(n6767), .C1(
        pipeline_regfile_data[697]), .C2(n6764), .A(n9075), .ZN(n9074) );
  OAI22_X2 U9472 ( .A1(n9076), .A2(n9305), .B1(n9077), .B2(n9306), .ZN(n9075)
         );
  NAND2_X2 U9473 ( .A1(n9081), .A2(n9082), .ZN(n9080) );
  NAND2_X2 U9474 ( .A1(pipeline_regfile_data[505]), .A2(n9320), .ZN(n9082) );
  NAND2_X2 U9475 ( .A1(pipeline_regfile_data[441]), .A2(n9321), .ZN(n9081) );
  AOI221_X2 U9476 ( .B1(pipeline_regfile_data[345]), .B2(n9323), .C1(
        pipeline_regfile_data[281]), .C2(n9326), .A(n9083), .ZN(n9078) );
  NAND2_X2 U9477 ( .A1(n9084), .A2(n9085), .ZN(n9083) );
  NAND2_X2 U9478 ( .A1(pipeline_regfile_data[473]), .A2(n9328), .ZN(n9085) );
  NAND2_X2 U9479 ( .A1(pipeline_regfile_data[409]), .A2(n9329), .ZN(n9084) );
  AND2_X1 U9480 ( .A1(n9086), .A2(n9087), .ZN(n9076) );
  NAND2_X2 U9481 ( .A1(n9089), .A2(n9090), .ZN(n9088) );
  NAND2_X2 U9482 ( .A1(pipeline_regfile_data[249]), .A2(n9320), .ZN(n9090) );
  NAND2_X2 U9483 ( .A1(pipeline_regfile_data[185]), .A2(n9321), .ZN(n9089) );
  AOI221_X2 U9484 ( .B1(pipeline_regfile_data[89]), .B2(n9323), .C1(
        pipeline_regfile_data[25]), .C2(n9327), .A(n9091), .ZN(n9086) );
  NAND2_X2 U9485 ( .A1(n9092), .A2(n9093), .ZN(n9091) );
  NAND2_X2 U9486 ( .A1(pipeline_regfile_data[217]), .A2(n9328), .ZN(n9093) );
  NAND2_X2 U9487 ( .A1(pipeline_regfile_data[153]), .A2(n9330), .ZN(n9092) );
  AOI221_X2 U9488 ( .B1(pipeline_regfile_data[1017]), .B2(n6765), .C1(
        pipeline_regfile_data[761]), .C2(n6761), .A(n9094), .ZN(n9073) );
  INV_X4 U9489 ( .A(n9095), .ZN(n9094) );
  AOI221_X2 U9490 ( .B1(pipeline_regfile_data[569]), .B2(n8299), .C1(
        pipeline_regfile_data[825]), .C2(n8300), .A(n9096), .ZN(n9095) );
  AND2_X1 U9491 ( .A1(pipeline_regfile_data[633]), .A2(n8302), .ZN(n9096) );
  NAND2_X2 U9492 ( .A1(n9098), .A2(n9099), .ZN(n9097) );
  NAND2_X2 U9493 ( .A1(pipeline_regfile_data[665]), .A2(n6769), .ZN(n9099) );
  NAND2_X2 U9494 ( .A1(pipeline_regfile_data[889]), .A2(n6770), .ZN(n9098) );
  AOI221_X2 U9495 ( .B1(pipeline_regfile_data[537]), .B2(n6709), .C1(
        pipeline_regfile_data[985]), .C2(n6763), .A(n9100), .ZN(n9071) );
  INV_X4 U9496 ( .A(n9101), .ZN(n9100) );
  AOI221_X2 U9497 ( .B1(pipeline_regfile_data[793]), .B2(n6766), .C1(
        pipeline_regfile_data[601]), .C2(n6762), .A(n9102), .ZN(n9101) );
  AND2_X1 U9498 ( .A1(pipeline_regfile_data[857]), .A2(n6768), .ZN(n9102) );
  AOI221_X2 U9499 ( .B1(pipeline_regfile_data[954]), .B2(n6767), .C1(
        pipeline_regfile_data[698]), .C2(n6764), .A(n9107), .ZN(n9106) );
  OAI22_X2 U9500 ( .A1(n9108), .A2(n9305), .B1(n9109), .B2(n9306), .ZN(n9107)
         );
  AND2_X1 U9501 ( .A1(n9110), .A2(n9111), .ZN(n9109) );
  AOI221_X2 U9502 ( .B1(pipeline_regfile_data[378]), .B2(n9308), .C1(
        pipeline_regfile_data[314]), .C2(n9313), .A(n9112), .ZN(n9111) );
  NAND2_X2 U9503 ( .A1(n9113), .A2(n9114), .ZN(n9112) );
  NAND2_X2 U9504 ( .A1(pipeline_regfile_data[506]), .A2(n9320), .ZN(n9114) );
  NAND2_X2 U9505 ( .A1(pipeline_regfile_data[442]), .A2(n9321), .ZN(n9113) );
  AOI221_X2 U9506 ( .B1(pipeline_regfile_data[346]), .B2(n9323), .C1(
        pipeline_regfile_data[282]), .C2(n9326), .A(n9115), .ZN(n9110) );
  NAND2_X2 U9507 ( .A1(n9116), .A2(n9117), .ZN(n9115) );
  NAND2_X2 U9508 ( .A1(pipeline_regfile_data[474]), .A2(n9328), .ZN(n9117) );
  NAND2_X2 U9509 ( .A1(pipeline_regfile_data[410]), .A2(n9329), .ZN(n9116) );
  AND2_X1 U9510 ( .A1(n9118), .A2(n9119), .ZN(n9108) );
  AOI221_X2 U9511 ( .B1(pipeline_regfile_data[122]), .B2(n9309), .C1(
        pipeline_regfile_data[58]), .C2(n9313), .A(n9120), .ZN(n9119) );
  NAND2_X2 U9512 ( .A1(n9121), .A2(n9122), .ZN(n9120) );
  NAND2_X2 U9513 ( .A1(pipeline_regfile_data[250]), .A2(n9318), .ZN(n9122) );
  NAND2_X2 U9514 ( .A1(pipeline_regfile_data[186]), .A2(n9321), .ZN(n9121) );
  NAND2_X2 U9515 ( .A1(n9124), .A2(n9125), .ZN(n9123) );
  NAND2_X2 U9516 ( .A1(pipeline_regfile_data[218]), .A2(n9328), .ZN(n9125) );
  NAND2_X2 U9517 ( .A1(pipeline_regfile_data[154]), .A2(n9330), .ZN(n9124) );
  AOI221_X2 U9518 ( .B1(pipeline_regfile_data[1018]), .B2(n6765), .C1(
        pipeline_regfile_data[762]), .C2(n6761), .A(n9126), .ZN(n9105) );
  INV_X4 U9519 ( .A(n9127), .ZN(n9126) );
  AOI221_X2 U9520 ( .B1(pipeline_regfile_data[570]), .B2(n8299), .C1(
        pipeline_regfile_data[826]), .C2(n8300), .A(n9128), .ZN(n9127) );
  AND2_X1 U9521 ( .A1(pipeline_regfile_data[634]), .A2(n8302), .ZN(n9128) );
  NAND2_X2 U9522 ( .A1(n9130), .A2(n9131), .ZN(n9129) );
  NAND2_X2 U9523 ( .A1(pipeline_regfile_data[666]), .A2(n6769), .ZN(n9131) );
  NAND2_X2 U9524 ( .A1(pipeline_regfile_data[890]), .A2(n6770), .ZN(n9130) );
  AOI221_X2 U9525 ( .B1(pipeline_regfile_data[538]), .B2(n6709), .C1(
        pipeline_regfile_data[986]), .C2(n6763), .A(n9132), .ZN(n9103) );
  INV_X4 U9526 ( .A(n9133), .ZN(n9132) );
  AOI221_X2 U9527 ( .B1(pipeline_regfile_data[794]), .B2(n6766), .C1(
        pipeline_regfile_data[602]), .C2(n6762), .A(n9134), .ZN(n9133) );
  AND2_X1 U9528 ( .A1(pipeline_regfile_data[858]), .A2(n6768), .ZN(n9134) );
  AOI221_X2 U9529 ( .B1(pipeline_regfile_data[955]), .B2(n6767), .C1(
        pipeline_regfile_data[699]), .C2(n6764), .A(n9139), .ZN(n9138) );
  OAI22_X2 U9530 ( .A1(n9140), .A2(n9305), .B1(n9141), .B2(n9306), .ZN(n9139)
         );
  AOI221_X2 U9531 ( .B1(pipeline_regfile_data[379]), .B2(n9308), .C1(
        pipeline_regfile_data[315]), .C2(n9313), .A(n9144), .ZN(n9143) );
  NAND2_X2 U9532 ( .A1(n9145), .A2(n9146), .ZN(n9144) );
  NAND2_X2 U9533 ( .A1(pipeline_regfile_data[507]), .A2(n9320), .ZN(n9146) );
  NAND2_X2 U9534 ( .A1(pipeline_regfile_data[443]), .A2(n9321), .ZN(n9145) );
  AOI221_X2 U9535 ( .B1(pipeline_regfile_data[347]), .B2(n9323), .C1(
        pipeline_regfile_data[283]), .C2(n9326), .A(n9147), .ZN(n9142) );
  NAND2_X2 U9536 ( .A1(n9148), .A2(n9149), .ZN(n9147) );
  NAND2_X2 U9537 ( .A1(pipeline_regfile_data[475]), .A2(n9328), .ZN(n9149) );
  NAND2_X2 U9538 ( .A1(pipeline_regfile_data[411]), .A2(n9329), .ZN(n9148) );
  AND2_X1 U9539 ( .A1(n9150), .A2(n9151), .ZN(n9140) );
  AOI221_X2 U9540 ( .B1(pipeline_regfile_data[123]), .B2(n9308), .C1(
        pipeline_regfile_data[59]), .C2(n9313), .A(n9152), .ZN(n9151) );
  NAND2_X2 U9541 ( .A1(n9153), .A2(n9154), .ZN(n9152) );
  NAND2_X2 U9542 ( .A1(pipeline_regfile_data[251]), .A2(n9319), .ZN(n9154) );
  NAND2_X2 U9543 ( .A1(pipeline_regfile_data[187]), .A2(n9321), .ZN(n9153) );
  AOI221_X2 U9544 ( .B1(pipeline_regfile_data[91]), .B2(n9323), .C1(
        pipeline_regfile_data[27]), .C2(n9326), .A(n9155), .ZN(n9150) );
  NAND2_X2 U9545 ( .A1(n9156), .A2(n9157), .ZN(n9155) );
  NAND2_X2 U9546 ( .A1(pipeline_regfile_data[219]), .A2(n9328), .ZN(n9157) );
  NAND2_X2 U9547 ( .A1(pipeline_regfile_data[155]), .A2(n9332), .ZN(n9156) );
  AOI221_X2 U9548 ( .B1(pipeline_regfile_data[1019]), .B2(n6765), .C1(
        pipeline_regfile_data[763]), .C2(n6761), .A(n9158), .ZN(n9137) );
  INV_X4 U9549 ( .A(n9159), .ZN(n9158) );
  AOI221_X2 U9550 ( .B1(pipeline_regfile_data[571]), .B2(n8299), .C1(
        pipeline_regfile_data[827]), .C2(n8300), .A(n9160), .ZN(n9159) );
  AND2_X1 U9551 ( .A1(pipeline_regfile_data[635]), .A2(n8302), .ZN(n9160) );
  AOI221_X2 U9552 ( .B1(pipeline_regfile_data[731]), .B2(n6773), .C1(
        pipeline_regfile_data[923]), .C2(n6772), .A(n9161), .ZN(n9136) );
  NAND2_X2 U9553 ( .A1(n9162), .A2(n9163), .ZN(n9161) );
  NAND2_X2 U9554 ( .A1(pipeline_regfile_data[667]), .A2(n6769), .ZN(n9163) );
  NAND2_X2 U9555 ( .A1(pipeline_regfile_data[891]), .A2(n6770), .ZN(n9162) );
  AOI221_X2 U9556 ( .B1(pipeline_regfile_data[539]), .B2(n6709), .C1(
        pipeline_regfile_data[987]), .C2(n6763), .A(n9164), .ZN(n9135) );
  INV_X4 U9557 ( .A(n9165), .ZN(n9164) );
  AOI221_X2 U9558 ( .B1(pipeline_regfile_data[795]), .B2(n6766), .C1(
        pipeline_regfile_data[603]), .C2(n6762), .A(n9166), .ZN(n9165) );
  AND2_X1 U9559 ( .A1(pipeline_regfile_data[859]), .A2(n6768), .ZN(n9166) );
  AOI221_X2 U9560 ( .B1(pipeline_regfile_data[956]), .B2(n6767), .C1(
        pipeline_regfile_data[700]), .C2(n6764), .A(n9171), .ZN(n9170) );
  OAI22_X2 U9561 ( .A1(n9172), .A2(n9305), .B1(n9173), .B2(n9306), .ZN(n9171)
         );
  AND2_X1 U9562 ( .A1(n9174), .A2(n9175), .ZN(n9173) );
  AOI221_X2 U9563 ( .B1(pipeline_regfile_data[380]), .B2(n9308), .C1(
        pipeline_regfile_data[316]), .C2(n9313), .A(n9176), .ZN(n9175) );
  NAND2_X2 U9564 ( .A1(n9177), .A2(n9178), .ZN(n9176) );
  NAND2_X2 U9565 ( .A1(pipeline_regfile_data[508]), .A2(n9319), .ZN(n9178) );
  NAND2_X2 U9566 ( .A1(pipeline_regfile_data[444]), .A2(n9321), .ZN(n9177) );
  AOI221_X2 U9567 ( .B1(pipeline_regfile_data[348]), .B2(n9323), .C1(
        pipeline_regfile_data[284]), .C2(n9326), .A(n9179), .ZN(n9174) );
  NAND2_X2 U9568 ( .A1(n9180), .A2(n9181), .ZN(n9179) );
  NAND2_X2 U9569 ( .A1(pipeline_regfile_data[476]), .A2(n9328), .ZN(n9181) );
  NAND2_X2 U9570 ( .A1(pipeline_regfile_data[412]), .A2(n9332), .ZN(n9180) );
  AND2_X1 U9571 ( .A1(n9182), .A2(n9183), .ZN(n9172) );
  AOI221_X2 U9572 ( .B1(pipeline_regfile_data[124]), .B2(n9308), .C1(
        pipeline_regfile_data[60]), .C2(n9313), .A(n9184), .ZN(n9183) );
  NAND2_X2 U9573 ( .A1(n9185), .A2(n9186), .ZN(n9184) );
  NAND2_X2 U9574 ( .A1(pipeline_regfile_data[252]), .A2(n9318), .ZN(n9186) );
  NAND2_X2 U9575 ( .A1(pipeline_regfile_data[188]), .A2(n9321), .ZN(n9185) );
  AOI221_X2 U9576 ( .B1(pipeline_regfile_data[92]), .B2(n9324), .C1(
        pipeline_regfile_data[28]), .C2(n9326), .A(n9187), .ZN(n9182) );
  NAND2_X2 U9577 ( .A1(n9188), .A2(n9189), .ZN(n9187) );
  NAND2_X2 U9578 ( .A1(pipeline_regfile_data[220]), .A2(n9328), .ZN(n9189) );
  NAND2_X2 U9579 ( .A1(pipeline_regfile_data[156]), .A2(n9330), .ZN(n9188) );
  AOI221_X2 U9580 ( .B1(pipeline_regfile_data[1020]), .B2(n6765), .C1(
        pipeline_regfile_data[764]), .C2(n6761), .A(n9190), .ZN(n9169) );
  INV_X4 U9581 ( .A(n9191), .ZN(n9190) );
  AOI221_X2 U9582 ( .B1(pipeline_regfile_data[572]), .B2(n8299), .C1(
        pipeline_regfile_data[828]), .C2(n8300), .A(n9192), .ZN(n9191) );
  AND2_X1 U9583 ( .A1(pipeline_regfile_data[636]), .A2(n8302), .ZN(n9192) );
  NAND2_X2 U9584 ( .A1(n9194), .A2(n9195), .ZN(n9193) );
  NAND2_X2 U9585 ( .A1(pipeline_regfile_data[668]), .A2(n6769), .ZN(n9195) );
  NAND2_X2 U9586 ( .A1(pipeline_regfile_data[892]), .A2(n6770), .ZN(n9194) );
  AOI221_X2 U9587 ( .B1(pipeline_regfile_data[540]), .B2(n6709), .C1(
        pipeline_regfile_data[988]), .C2(n6763), .A(n9196), .ZN(n9167) );
  INV_X4 U9588 ( .A(n9197), .ZN(n9196) );
  AOI221_X2 U9589 ( .B1(pipeline_regfile_data[796]), .B2(n6766), .C1(
        pipeline_regfile_data[604]), .C2(n6762), .A(n9198), .ZN(n9197) );
  AND2_X1 U9590 ( .A1(pipeline_regfile_data[860]), .A2(n6768), .ZN(n9198) );
  AOI221_X2 U9591 ( .B1(pipeline_regfile_data[957]), .B2(n6767), .C1(
        pipeline_regfile_data[701]), .C2(n6764), .A(n9203), .ZN(n9202) );
  OAI22_X2 U9592 ( .A1(n9204), .A2(n9305), .B1(n9205), .B2(n9306), .ZN(n9203)
         );
  AND2_X1 U9593 ( .A1(n9206), .A2(n9207), .ZN(n9205) );
  AOI221_X2 U9594 ( .B1(pipeline_regfile_data[381]), .B2(n9308), .C1(
        pipeline_regfile_data[317]), .C2(n9313), .A(n9208), .ZN(n9207) );
  NAND2_X2 U9595 ( .A1(n9209), .A2(n9210), .ZN(n9208) );
  NAND2_X2 U9596 ( .A1(pipeline_regfile_data[509]), .A2(n9320), .ZN(n9210) );
  NAND2_X2 U9597 ( .A1(pipeline_regfile_data[445]), .A2(n9321), .ZN(n9209) );
  AOI221_X2 U9598 ( .B1(pipeline_regfile_data[349]), .B2(n9323), .C1(
        pipeline_regfile_data[285]), .C2(n9327), .A(n9211), .ZN(n9206) );
  NAND2_X2 U9599 ( .A1(n9212), .A2(n9213), .ZN(n9211) );
  NAND2_X2 U9600 ( .A1(pipeline_regfile_data[477]), .A2(n9328), .ZN(n9213) );
  NAND2_X2 U9601 ( .A1(pipeline_regfile_data[413]), .A2(n9332), .ZN(n9212) );
  AND2_X1 U9602 ( .A1(n9214), .A2(n9215), .ZN(n9204) );
  AOI221_X2 U9603 ( .B1(pipeline_regfile_data[125]), .B2(n9308), .C1(
        pipeline_regfile_data[61]), .C2(n9313), .A(n9216), .ZN(n9215) );
  NAND2_X2 U9604 ( .A1(n9217), .A2(n9218), .ZN(n9216) );
  NAND2_X2 U9605 ( .A1(pipeline_regfile_data[253]), .A2(n9320), .ZN(n9218) );
  NAND2_X2 U9606 ( .A1(pipeline_regfile_data[189]), .A2(n9321), .ZN(n9217) );
  AOI221_X2 U9607 ( .B1(pipeline_regfile_data[93]), .B2(n9323), .C1(
        pipeline_regfile_data[29]), .C2(n9326), .A(n9219), .ZN(n9214) );
  NAND2_X2 U9608 ( .A1(n9220), .A2(n9221), .ZN(n9219) );
  NAND2_X2 U9609 ( .A1(pipeline_regfile_data[221]), .A2(n9328), .ZN(n9221) );
  NAND2_X2 U9610 ( .A1(pipeline_regfile_data[157]), .A2(n9329), .ZN(n9220) );
  AOI221_X2 U9611 ( .B1(pipeline_regfile_data[1021]), .B2(n6765), .C1(
        pipeline_regfile_data[765]), .C2(n6761), .A(n9222), .ZN(n9201) );
  INV_X4 U9612 ( .A(n9223), .ZN(n9222) );
  AOI221_X2 U9613 ( .B1(pipeline_regfile_data[573]), .B2(n8299), .C1(
        pipeline_regfile_data[829]), .C2(n8300), .A(n9224), .ZN(n9223) );
  AND2_X1 U9614 ( .A1(pipeline_regfile_data[637]), .A2(n8302), .ZN(n9224) );
  NAND2_X2 U9615 ( .A1(n9226), .A2(n9227), .ZN(n9225) );
  NAND2_X2 U9616 ( .A1(pipeline_regfile_data[669]), .A2(n6769), .ZN(n9227) );
  NAND2_X2 U9617 ( .A1(pipeline_regfile_data[893]), .A2(n6770), .ZN(n9226) );
  AOI221_X2 U9618 ( .B1(pipeline_regfile_data[541]), .B2(n6709), .C1(
        pipeline_regfile_data[989]), .C2(n6763), .A(n9228), .ZN(n9199) );
  INV_X4 U9619 ( .A(n9229), .ZN(n9228) );
  AOI221_X2 U9620 ( .B1(pipeline_regfile_data[797]), .B2(n6766), .C1(
        pipeline_regfile_data[605]), .C2(n6762), .A(n9230), .ZN(n9229) );
  AND2_X1 U9621 ( .A1(pipeline_regfile_data[861]), .A2(n6768), .ZN(n9230) );
  AOI221_X2 U9622 ( .B1(pipeline_regfile_data[958]), .B2(n6767), .C1(
        pipeline_regfile_data[702]), .C2(n6764), .A(n9235), .ZN(n9234) );
  OAI22_X2 U9623 ( .A1(n9236), .A2(n9305), .B1(n9237), .B2(n9306), .ZN(n9235)
         );
  AND2_X1 U9624 ( .A1(n9238), .A2(n9239), .ZN(n9237) );
  AOI221_X2 U9625 ( .B1(pipeline_regfile_data[382]), .B2(n9308), .C1(
        pipeline_regfile_data[318]), .C2(n9313), .A(n9240), .ZN(n9239) );
  NAND2_X2 U9626 ( .A1(n9241), .A2(n9242), .ZN(n9240) );
  NAND2_X2 U9627 ( .A1(pipeline_regfile_data[510]), .A2(n9319), .ZN(n9242) );
  NAND2_X2 U9628 ( .A1(pipeline_regfile_data[446]), .A2(n9321), .ZN(n9241) );
  AOI221_X2 U9629 ( .B1(pipeline_regfile_data[350]), .B2(n9323), .C1(
        pipeline_regfile_data[286]), .C2(n9326), .A(n9243), .ZN(n9238) );
  NAND2_X2 U9630 ( .A1(n9244), .A2(n9245), .ZN(n9243) );
  NAND2_X2 U9631 ( .A1(pipeline_regfile_data[478]), .A2(n9328), .ZN(n9245) );
  NAND2_X2 U9632 ( .A1(pipeline_regfile_data[414]), .A2(n9329), .ZN(n9244) );
  AND2_X1 U9633 ( .A1(n9246), .A2(n9247), .ZN(n9236) );
  AOI221_X2 U9634 ( .B1(pipeline_regfile_data[126]), .B2(n9308), .C1(
        pipeline_regfile_data[62]), .C2(n9313), .A(n9248), .ZN(n9247) );
  NAND2_X2 U9635 ( .A1(n9249), .A2(n9250), .ZN(n9248) );
  NAND2_X2 U9636 ( .A1(pipeline_regfile_data[254]), .A2(n9318), .ZN(n9250) );
  NAND2_X2 U9637 ( .A1(pipeline_regfile_data[190]), .A2(n9321), .ZN(n9249) );
  AOI221_X2 U9638 ( .B1(pipeline_regfile_data[94]), .B2(n9324), .C1(
        pipeline_regfile_data[30]), .C2(n9326), .A(n9251), .ZN(n9246) );
  NAND2_X2 U9639 ( .A1(n9252), .A2(n9253), .ZN(n9251) );
  NAND2_X2 U9640 ( .A1(pipeline_regfile_data[222]), .A2(n9328), .ZN(n9253) );
  NAND2_X2 U9641 ( .A1(pipeline_regfile_data[158]), .A2(n9330), .ZN(n9252) );
  AOI221_X2 U9642 ( .B1(pipeline_regfile_data[1022]), .B2(n6765), .C1(
        pipeline_regfile_data[766]), .C2(n6761), .A(n9254), .ZN(n9233) );
  INV_X4 U9643 ( .A(n9255), .ZN(n9254) );
  AOI221_X2 U9644 ( .B1(pipeline_regfile_data[574]), .B2(n8299), .C1(
        pipeline_regfile_data[830]), .C2(n8300), .A(n9256), .ZN(n9255) );
  AND2_X1 U9645 ( .A1(pipeline_regfile_data[638]), .A2(n8302), .ZN(n9256) );
  NAND2_X2 U9646 ( .A1(n9258), .A2(n9259), .ZN(n9257) );
  NAND2_X2 U9647 ( .A1(pipeline_regfile_data[670]), .A2(n6769), .ZN(n9259) );
  NAND2_X2 U9648 ( .A1(pipeline_regfile_data[894]), .A2(n6770), .ZN(n9258) );
  AOI221_X2 U9649 ( .B1(pipeline_regfile_data[542]), .B2(n6709), .C1(
        pipeline_regfile_data[990]), .C2(n6763), .A(n9260), .ZN(n9231) );
  INV_X4 U9650 ( .A(n9261), .ZN(n9260) );
  AOI221_X2 U9651 ( .B1(pipeline_regfile_data[798]), .B2(n6766), .C1(
        pipeline_regfile_data[606]), .C2(n6762), .A(n9262), .ZN(n9261) );
  AND2_X1 U9652 ( .A1(pipeline_regfile_data[862]), .A2(n6768), .ZN(n9262) );
  OAI22_X2 U9653 ( .A1(n9268), .A2(n9305), .B1(n9269), .B2(n9306), .ZN(n9267)
         );
  AND2_X1 U9654 ( .A1(n9271), .A2(n9272), .ZN(n9269) );
  AOI221_X2 U9655 ( .B1(pipeline_regfile_data[383]), .B2(n9308), .C1(
        pipeline_regfile_data[319]), .C2(n9313), .A(n9273), .ZN(n9272) );
  NAND2_X2 U9656 ( .A1(n9274), .A2(n9275), .ZN(n9273) );
  NAND2_X2 U9657 ( .A1(pipeline_regfile_data[511]), .A2(n9320), .ZN(n9275) );
  NAND2_X2 U9658 ( .A1(pipeline_regfile_data[447]), .A2(n9321), .ZN(n9274) );
  AOI221_X2 U9659 ( .B1(pipeline_regfile_data[351]), .B2(n9323), .C1(
        pipeline_regfile_data[287]), .C2(n9327), .A(n9276), .ZN(n9271) );
  NAND2_X2 U9660 ( .A1(n9277), .A2(n9278), .ZN(n9276) );
  NAND2_X2 U9661 ( .A1(pipeline_regfile_data[479]), .A2(n9328), .ZN(n9278) );
  NAND2_X2 U9662 ( .A1(n9279), .A2(n9270), .ZN(n8278) );
  AND2_X1 U9663 ( .A1(n9280), .A2(n9281), .ZN(n9268) );
  AOI221_X2 U9664 ( .B1(pipeline_regfile_data[127]), .B2(n9308), .C1(
        pipeline_regfile_data[63]), .C2(n9313), .A(n9282), .ZN(n9281) );
  NAND2_X2 U9665 ( .A1(n9283), .A2(n9284), .ZN(n9282) );
  NAND2_X2 U9666 ( .A1(pipeline_regfile_data[255]), .A2(n9319), .ZN(n9284) );
  NAND2_X2 U9667 ( .A1(pipeline_regfile_data[191]), .A2(n9321), .ZN(n9283) );
  AOI221_X2 U9668 ( .B1(pipeline_regfile_data[95]), .B2(n9323), .C1(
        pipeline_regfile_data[31]), .C2(n9326), .A(n9285), .ZN(n9280) );
  NAND2_X2 U9669 ( .A1(n9286), .A2(n9287), .ZN(n9285) );
  NAND2_X2 U9670 ( .A1(pipeline_regfile_data[223]), .A2(n9328), .ZN(n9287) );
  NAND2_X2 U9671 ( .A1(pipeline_regfile_data[159]), .A2(n9330), .ZN(n9286) );
  AOI221_X2 U9672 ( .B1(pipeline_regfile_data[1023]), .B2(n6765), .C1(
        pipeline_regfile_data[767]), .C2(n6761), .A(n9288), .ZN(n9265) );
  INV_X4 U9673 ( .A(n9289), .ZN(n9288) );
  AOI221_X2 U9674 ( .B1(pipeline_regfile_data[575]), .B2(n8299), .C1(
        pipeline_regfile_data[831]), .C2(n8300), .A(n9290), .ZN(n9289) );
  AND2_X1 U9675 ( .A1(pipeline_regfile_data[639]), .A2(n8302), .ZN(n9290) );
  NAND2_X2 U9676 ( .A1(n9313), .A2(n7164), .ZN(n9292) );
  NAND2_X2 U9677 ( .A1(n9296), .A2(n9297), .ZN(n9295) );
  NAND2_X2 U9678 ( .A1(pipeline_regfile_data[671]), .A2(n6769), .ZN(n9297) );
  NAND2_X2 U9679 ( .A1(pipeline_regfile_data[895]), .A2(n6770), .ZN(n9296) );
  AOI221_X2 U9680 ( .B1(pipeline_regfile_data[543]), .B2(n6709), .C1(
        pipeline_regfile_data[991]), .C2(n6763), .A(n9299), .ZN(n9263) );
  INV_X4 U9681 ( .A(n9300), .ZN(n9299) );
  AOI221_X2 U9682 ( .B1(pipeline_regfile_data[799]), .B2(n6766), .C1(
        pipeline_regfile_data[607]), .C2(n6762), .A(n9301), .ZN(n9300) );
  AND2_X1 U9683 ( .A1(pipeline_regfile_data[863]), .A2(n6768), .ZN(n9301) );
  INV_X4 U9684 ( .A(n9302), .ZN(n8285) );
  NAND3_X1 U9685 ( .A1(pipeline_regfile_N14), .A2(pipeline_regfile_N13), .A3(
        n636), .ZN(n9303) );
  NAND3_X1 U9686 ( .A1(pipeline_regfile_N13), .A2(n638), .A3(n636), .ZN(n9302)
         );
  NAND2_X1 U9687 ( .A1(n12180), .A2(pipeline_alu_src_b[27]), .ZN(n12181) );
  NOR2_X1 U9688 ( .A1(pipeline_alu_src_b[27]), .A2(n12357), .ZN(n12166) );
  INV_X1 U9689 ( .A(pipeline_alu_src_b[27]), .ZN(n10027) );
  OAI221_X4 U9690 ( .B1(n10026), .B2(n9448), .C1(n10236), .C2(n9397), .A(
        n10043), .ZN(pipeline_alu_src_b[27]) );
  AOI221_X1 U9691 ( .B1(pipeline_regfile_N13), .B2(n10332), .C1(n6666), .C2(
        n6637), .A(n10331), .ZN(n1911) );
  XNOR2_X1 U9692 ( .A(pipeline_reg_to_wr_WB[1]), .B(pipeline_regfile_N13), 
        .ZN(n9647) );
  INV_X2 U9693 ( .A(n9391), .ZN(n9442) );
  INV_X4 U9694 ( .A(n13174), .ZN(n10808) );
  NAND2_X1 U9695 ( .A1(n9385), .A2(n9892), .ZN(n9896) );
  NAND4_X1 U9696 ( .A1(n12149), .A2(n13130), .A3(n12621), .A4(n12150), .ZN(
        n12620) );
  NAND3_X1 U9697 ( .A1(n12600), .A2(n12149), .A3(n12148), .ZN(n12150) );
  NOR2_X1 U9698 ( .A1(pipeline_rs1_data_bypassed[12]), .A2(n9463), .ZN(n10878)
         );
  AOI221_X1 U9699 ( .B1(pipeline_md_N41), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[12]), .A(n10854), .ZN(n10855) );
  OAI221_X1 U9700 ( .B1(n11280), .B2(n638), .C1(n12530), .C2(n9467), .A(n10415), .ZN(n10416) );
  OAI22_X1 U9701 ( .A1(n603), .A2(n637), .B1(n6636), .B2(pipeline_dmem_type_2_), .ZN(n10330) );
  NOR2_X1 U9702 ( .A1(pipeline_rs1_data_bypassed[11]), .A2(n9463), .ZN(n10932)
         );
  AOI221_X1 U9703 ( .B1(pipeline_md_N40), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[11]), .A(n10908), .ZN(n10909) );
  NAND3_X1 U9704 ( .A1(pipeline_regfile_N17), .A2(n7163), .A3(n6847), .ZN(
        n11323) );
  NAND3_X1 U9705 ( .A1(n6748), .A2(pipeline_regfile_N17), .A3(n7174), .ZN(
        n12806) );
  NAND2_X1 U9707 ( .A1(n9790), .A2(pipeline_regfile_N17), .ZN(n9719) );
  INV_X4 U9709 ( .A(pipeline_alu_src_a[8]), .ZN(n9334) );
  INV_X1 U9710 ( .A(n9334), .ZN(n9335) );
  OAI22_X1 U9711 ( .A1(n12274), .A2(n12565), .B1(n6619), .B2(n9400), .ZN(
        n12275) );
  NAND2_X1 U9712 ( .A1(n12411), .A2(n12560), .ZN(n12410) );
  NOR4_X1 U9713 ( .A1(n10080), .A2(n12398), .A3(n10079), .A4(n10078), .ZN(
        n10089) );
  NAND2_X2 U9714 ( .A1(n12561), .A2(n12557), .ZN(n9336) );
  NOR2_X1 U9715 ( .A1(ext_interrupts[8]), .A2(n6960), .ZN(n9591) );
  AOI22_X2 U9716 ( .A1(ext_interrupts[8]), .A2(n9564), .B1(ext_interrupts[7]), 
        .B2(n11114), .ZN(n9567) );
  INV_X1 U9717 ( .A(ext_interrupts[10]), .ZN(n13137) );
  NOR2_X1 U9718 ( .A1(ext_interrupts[11]), .A2(ext_interrupts[10]), .ZN(n9592)
         );
  AOI22_X2 U9719 ( .A1(ext_interrupts[11]), .A2(n9562), .B1(ext_interrupts[10]), .B2(pipeline_csr_mie[18]), .ZN(n9569) );
  INV_X2 U9720 ( .A(n9884), .ZN(n9872) );
  NAND3_X1 U9721 ( .A1(n793), .A2(n6369), .A3(n10348), .ZN(n10349) );
  NAND2_X1 U9723 ( .A1(n10348), .A2(n9676), .ZN(n12395) );
  AOI221_X1 U9724 ( .B1(pipeline_md_N34), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[5]), .A(n10769), .ZN(n10770) );
  NOR2_X1 U9725 ( .A1(pipeline_rs1_data_bypassed[5]), .A2(n9463), .ZN(n10791)
         );
  AOI221_X1 U9726 ( .B1(pipeline_md_N67), .B2(n6797), .C1(n12749), .C2(n7004), 
        .A(n12740), .ZN(n12741) );
  AOI221_X1 U9727 ( .B1(pipeline_md_N64), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[1]), .A(n12746), .ZN(n12747) );
  INV_X2 U9728 ( .A(n9871), .ZN(n9867) );
  AOI221_X1 U9729 ( .B1(pipeline_md_N35), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[6]), .A(n10718), .ZN(n10719) );
  NOR2_X1 U9730 ( .A1(pipeline_rs1_data_bypassed[6]), .A2(n9463), .ZN(n10739)
         );
  AOI221_X1 U9731 ( .B1(pipeline_md_N71), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[8]), .A(n12732), .ZN(n12733) );
  AOI221_X1 U9732 ( .B1(pipeline_md_N31), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[2]), .A(n10390), .ZN(n10391) );
  AOI221_X1 U9733 ( .B1(n603), .B2(pipeline_rs1_data_bypassed[2]), .C1(
        pipeline_regfile_N14), .C2(pipeline_dmem_type_2_), .A(n10413), .ZN(
        n10414) );
  INV_X4 U9734 ( .A(n13185), .ZN(n9340) );
  INV_X4 U9735 ( .A(n13183), .ZN(n9342) );
  INV_X4 U9736 ( .A(n13184), .ZN(n9344) );
  INV_X4 U9737 ( .A(n13175), .ZN(n9346) );
  INV_X4 U9738 ( .A(n13176), .ZN(n9348) );
  INV_X4 U9739 ( .A(n13177), .ZN(n9350) );
  INV_X4 U9740 ( .A(n13178), .ZN(n9352) );
  INV_X4 U9741 ( .A(n13179), .ZN(n9354) );
  INV_X4 U9742 ( .A(n13180), .ZN(n9356) );
  INV_X4 U9743 ( .A(n13181), .ZN(n9358) );
  INV_X4 U9744 ( .A(n13172), .ZN(n9362) );
  INV_X4 U9745 ( .A(n13166), .ZN(n9364) );
  INV_X4 U9746 ( .A(n13169), .ZN(n9366) );
  INV_X4 U9747 ( .A(n13171), .ZN(n9368) );
  INV_X4 U9748 ( .A(n13173), .ZN(n9374) );
  INV_X4 U9749 ( .A(n13170), .ZN(n9376) );
  INV_X4 U9750 ( .A(n13164), .ZN(n9378) );
  AOI221_X1 U9751 ( .B1(pipeline_md_N75), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[12]), .A(n12724), .ZN(n12725) );
  INV_X4 U9752 ( .A(pipeline_alu_src_b[4]), .ZN(n12800) );
  AND2_X4 U9753 ( .A1(n7178), .A2(n9723), .ZN(n9386) );
  OAI22_X1 U9754 ( .A1(n12792), .A2(n12565), .B1(n6610), .B2(n9401), .ZN(n9783) );
  AOI221_X1 U9755 ( .B1(n9471), .B2(n6619), .C1(n12276), .C2(n12792), .A(
        n11165), .ZN(n11755) );
  AOI221_X1 U9756 ( .B1(pipeline_md_N39), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[10]), .A(n10962), .ZN(n10963) );
  NOR2_X1 U9757 ( .A1(pipeline_rs1_data_bypassed[10]), .A2(n9463), .ZN(n10986)
         );
  AOI221_X1 U9758 ( .B1(n11506), .B2(n6571), .C1(n12062), .C2(n12094), .A(
        n11505), .ZN(n11516) );
  NAND2_X1 U9759 ( .A1(n9471), .A2(n6572), .ZN(n11721) );
  NAND2_X1 U9760 ( .A1(n11869), .A2(n6572), .ZN(n11871) );
  OAI22_X1 U9761 ( .A1(n6572), .A2(n12565), .B1(n6612), .B2(n9400), .ZN(n11169) );
  OAI22_X1 U9762 ( .A1(n6567), .A2(n12565), .B1(n6571), .B2(n12273), .ZN(
        n11401) );
  AOI221_X1 U9763 ( .B1(n9471), .B2(n6973), .C1(n12276), .C2(n6571), .A(n9762), 
        .ZN(n12775) );
  INV_X2 U9764 ( .A(n9925), .ZN(n9917) );
  AOI221_X1 U9765 ( .B1(n11649), .B2(pipeline_alu_src_a[12]), .C1(n12062), 
        .C2(n12226), .A(n11648), .ZN(n11659) );
  AOI221_X1 U9766 ( .B1(n9471), .B2(n11573), .C1(n12276), .C2(n6924), .A(
        n11168), .ZN(n11758) );
  OAI221_X1 U9767 ( .B1(n6924), .B2(n11574), .C1(n11573), .C2(n11572), .A(
        n11571), .ZN(n12135) );
  NAND2_X1 U9768 ( .A1(n11869), .A2(pipeline_alu_src_a[12]), .ZN(n11720) );
  AOI221_X1 U9769 ( .B1(n9471), .B2(n6924), .C1(n12276), .C2(n6613), .A(n11401), .ZN(n11675) );
  OAI22_X1 U9770 ( .A1(pipeline_alu_src_a[12]), .A2(n12565), .B1(n6973), .B2(
        n9401), .ZN(n11367) );
  AOI221_X1 U9771 ( .B1(n9471), .B2(n6614), .C1(n12276), .C2(
        pipeline_alu_src_a[12]), .A(n11497), .ZN(n12278) );
  OAI22_X1 U9772 ( .A1(n6924), .A2(n12565), .B1(n11414), .B2(n9400), .ZN(n9771) );
  AOI221_X1 U9773 ( .B1(n12363), .B2(n12362), .C1(n12361), .C2(n6976), .A(
        n12360), .ZN(n12381) );
  NOR2_X1 U9774 ( .A1(n6976), .A2(n12357), .ZN(n12358) );
  NAND2_X1 U9775 ( .A1(n7005), .A2(n6976), .ZN(n11411) );
  NAND2_X1 U9776 ( .A1(n6976), .A2(n6617), .ZN(n9400) );
  NAND2_X1 U9777 ( .A1(n6976), .A2(n6618), .ZN(n12273) );
  NAND2_X1 U9778 ( .A1(n6976), .A2(n11404), .ZN(n11572) );
  NAND2_X1 U9779 ( .A1(n6976), .A2(n6617), .ZN(n9401) );
  INV_X2 U9780 ( .A(n9869), .ZN(n9870) );
  AOI221_X1 U9781 ( .B1(pipeline_md_N70), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[7]), .A(n12734), .ZN(n12735) );
  NAND2_X1 U9782 ( .A1(n9848), .A2(n9849), .ZN(n9853) );
  INV_X2 U9783 ( .A(n9849), .ZN(n9851) );
  INV_X4 U9784 ( .A(pipeline_alu_src_b[8]), .ZN(n9387) );
  INV_X8 U9785 ( .A(n9483), .ZN(n9484) );
  OAI21_X2 U9786 ( .B1(n9901), .B2(n9845), .A(n9900), .ZN(n9906) );
  OAI21_X2 U9787 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9905) );
  AND2_X1 U9788 ( .A1(n7178), .A2(n9723), .ZN(n9390) );
  INV_X4 U9789 ( .A(n9657), .ZN(n9389) );
  AND2_X4 U9790 ( .A1(n9389), .A2(n7178), .ZN(n9724) );
  OAI22_X1 U9791 ( .A1(pipeline_alu_src_a[18]), .A2(n12565), .B1(n6597), .B2(
        n12273), .ZN(n11473) );
  OAI22_X1 U9792 ( .A1(n6598), .A2(n12565), .B1(pipeline_alu_src_a[12]), .B2(
        n9401), .ZN(n11343) );
  AOI221_X1 U9793 ( .B1(n9471), .B2(pipeline_alu_src_a[14]), .C1(n12276), .C2(
        n6597), .A(n11436), .ZN(n12371) );
  INV_X4 U9794 ( .A(n6596), .ZN(n11414) );
  AOI221_X1 U9795 ( .B1(pipeline_md_N45), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[16]), .A(n11069), .ZN(n11070) );
  NOR2_X1 U9796 ( .A1(pipeline_rs1_data_bypassed[16]), .A2(n9463), .ZN(n11093)
         );
  OAI22_X1 U9797 ( .A1(pipeline_alu_src_a[16]), .A2(n12565), .B1(n6567), .B2(
        n9401), .ZN(n11377) );
  OAI22_X1 U9798 ( .A1(pipeline_alu_src_a[19]), .A2(n12565), .B1(
        pipeline_alu_src_a[16]), .B2(n9401), .ZN(n11545) );
  NAND2_X1 U9799 ( .A1(n9489), .A2(pipeline_alu_src_a[16]), .ZN(n9747) );
  AOI221_X1 U9800 ( .B1(n11806), .B2(n6605), .C1(n12062), .C2(n11805), .A(
        n11804), .ZN(n11813) );
  OAI22_X1 U9801 ( .A1(n6606), .A2(n12565), .B1(n6635), .B2(n9400), .ZN(n11165) );
  NAND2_X1 U9802 ( .A1(n11869), .A2(n6606), .ZN(n12130) );
  NAND2_X1 U9803 ( .A1(n9471), .A2(n6605), .ZN(n11717) );
  AOI221_X1 U9804 ( .B1(n9471), .B2(n6621), .C1(n12276), .C2(n6606), .A(n9783), 
        .ZN(n12777) );
  INV_X2 U9805 ( .A(n9899), .ZN(n9845) );
  INV_X4 U9806 ( .A(n9442), .ZN(n9441) );
  AOI221_X1 U9807 ( .B1(pipeline_md_N37), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[8]), .A(n10610), .ZN(n10611) );
  NOR2_X1 U9808 ( .A1(pipeline_rs1_data_bypassed[8]), .A2(n9463), .ZN(n10632)
         );
  AOI221_X1 U9809 ( .B1(n11990), .B2(n9335), .C1(n12062), .C2(n11989), .A(
        n11988), .ZN(n11996) );
  AOI221_X1 U9810 ( .B1(n9471), .B2(n6612), .C1(n12276), .C2(n9335), .A(n11799), .ZN(n12272) );
  OAI22_X1 U9811 ( .A1(n9335), .A2(n12565), .B1(n6620), .B2(n9400), .ZN(n11368) );
  NAND2_X1 U9812 ( .A1(n9471), .A2(n9335), .ZN(n11873) );
  NAND2_X1 U9813 ( .A1(n11869), .A2(n9335), .ZN(n11715) );
  NAND2_X1 U9814 ( .A1(n12600), .A2(n12599), .ZN(n12624) );
  NOR2_X1 U9815 ( .A1(n6633), .A2(n12123), .ZN(n12124) );
  AOI221_X1 U9816 ( .B1(n9471), .B2(n6633), .C1(n12276), .C2(n12274), .A(
        n11365), .ZN(n11366) );
  OAI221_X1 U9817 ( .B1(n12274), .B2(n11572), .C1(n6633), .C2(n9401), .A(n9772), .ZN(n9773) );
  INV_X2 U9818 ( .A(n9868), .ZN(n9394) );
  NOR2_X2 U9819 ( .A1(n9597), .A2(n9598), .ZN(n9395) );
  NOR2_X1 U9820 ( .A1(n6631), .A2(n12359), .ZN(n12360) );
  NOR2_X1 U9821 ( .A1(n6575), .A2(n9724), .ZN(n9674) );
  AOI221_X1 U9822 ( .B1(pipeline_md_N33), .B2(n6798), .C1(n6808), .C2(n6998), 
        .A(n12675), .ZN(n12676) );
  NAND2_X1 U9823 ( .A1(n603), .A2(n6998), .ZN(n11245) );
  OAI21_X4 U9824 ( .B1(n10069), .B2(n10068), .A(n10067), .ZN(n12398) );
  AOI221_X1 U9825 ( .B1(pipeline_md_N66), .B2(n6797), .C1(n12749), .C2(n6987), 
        .A(n12742), .ZN(n12743) );
  AOI221_X1 U9826 ( .B1(n12363), .B2(n12126), .C1(n12125), .C2(n9339), .A(
        n12124), .ZN(n12142) );
  NOR2_X1 U9827 ( .A1(n9339), .A2(n12058), .ZN(n11584) );
  NOR3_X1 U9828 ( .A1(n12786), .A2(n9339), .A3(n12785), .ZN(n12787) );
  NOR2_X1 U9829 ( .A1(n9339), .A2(n12357), .ZN(n12122) );
  NAND2_X1 U9830 ( .A1(n7006), .A2(n9339), .ZN(n12027) );
  NAND2_X1 U9832 ( .A1(n9339), .A2(n9399), .ZN(n12645) );
  NAND3_X4 U9833 ( .A1(n12408), .A2(n12409), .A3(n12412), .ZN(n12557) );
  NAND3_X4 U9834 ( .A1(n12411), .A2(n12407), .A3(n12409), .ZN(n12561) );
  OAI221_X4 U9835 ( .B1(n598), .B2(n9795), .C1(n9792), .C2(n9448), .A(n9791), 
        .ZN(pipeline_alu_src_b[4]) );
  NAND2_X2 U9836 ( .A1(n9721), .A2(n12834), .ZN(n9396) );
  NAND2_X2 U9837 ( .A1(n9721), .A2(n12834), .ZN(n9397) );
  OAI22_X4 U9838 ( .A1(n744), .A2(n9445), .B1(n12422), .B2(n9443), .ZN(
        pipeline_alu_src_a[29]) );
  OAI22_X4 U9839 ( .A1(n733), .A2(n9445), .B1(n12466), .B2(n9443), .ZN(
        pipeline_alu_src_a[18]) );
  OAI22_X4 U9840 ( .A1(n729), .A2(n9445), .B1(n12481), .B2(n9443), .ZN(
        pipeline_alu_src_a[14]) );
  OAI221_X2 U9841 ( .B1(n12925), .B2(n12924), .C1(n12923), .C2(n9407), .A(
        n9411), .ZN(n9424) );
  OAI221_X2 U9842 ( .B1(n12925), .B2(n12924), .C1(n12923), .C2(n9407), .A(
        n9410), .ZN(n9425) );
  OAI221_X2 U9843 ( .B1(n12930), .B2(n12929), .C1(n12928), .C2(n9407), .A(
        n9410), .ZN(n9426) );
  OAI221_X2 U9844 ( .B1(n12930), .B2(n12929), .C1(n12928), .C2(n9407), .A(
        n12940), .ZN(n9427) );
  OAI221_X2 U9845 ( .B1(n12935), .B2(n12934), .C1(n12933), .C2(n9407), .A(
        n12940), .ZN(n9428) );
  OAI221_X2 U9846 ( .B1(n12935), .B2(n12934), .C1(n12933), .C2(n9407), .A(
        n9411), .ZN(n9429) );
  OAI221_X2 U9847 ( .B1(n12943), .B2(n12942), .C1(n12941), .C2(n9407), .A(
        n9411), .ZN(n9430) );
  OAI221_X2 U9848 ( .B1(n12943), .B2(n12942), .C1(n12941), .C2(n9407), .A(
        n9410), .ZN(n9431) );
  OAI22_X2 U9849 ( .A1(n12952), .A2(n9407), .B1(n12951), .B2(n12985), .ZN(
        n9432) );
  OAI22_X2 U9850 ( .A1(n12957), .A2(n9407), .B1(n12956), .B2(n12985), .ZN(
        n9433) );
  OAI22_X2 U9851 ( .A1(n12962), .A2(n9407), .B1(n12961), .B2(n12985), .ZN(
        n9434) );
  OAI22_X2 U9852 ( .A1(n12967), .A2(n9407), .B1(n12966), .B2(n12985), .ZN(
        n9435) );
  OAI22_X2 U9853 ( .A1(n12972), .A2(n9407), .B1(n12971), .B2(n12985), .ZN(
        n9436) );
  OAI22_X2 U9854 ( .A1(n12977), .A2(n9407), .B1(n12976), .B2(n12985), .ZN(
        n9437) );
  OAI22_X2 U9855 ( .A1(n12987), .A2(n9407), .B1(n12986), .B2(n12985), .ZN(
        n9438) );
  OR2_X1 U9856 ( .A1(dmem_hresp), .A2(pipeline_ctrl_had_ex_WB), .ZN(n12148)
         );
  INV_X4 U9857 ( .A(n12148), .ZN(n6369) );
  NAND2_X2 U9858 ( .A1(pipeline_csr_mie[8]), .A2(ext_interrupts[0]), .ZN(n9540) );
  NAND2_X2 U9859 ( .A1(ext_interrupts[1]), .A2(n9536), .ZN(n9539) );
  NAND2_X2 U9860 ( .A1(ext_interrupts[15]), .A2(n9537), .ZN(n9538) );
  NAND3_X2 U9861 ( .A1(n9540), .A2(n9539), .A3(n9538), .ZN(n9546) );
  NAND2_X2 U9862 ( .A1(pipeline_csr_mie[10]), .A2(ext_interrupts[2]), .ZN(
        n9544) );
  NAND2_X2 U9863 ( .A1(pipeline_csr_mie[11]), .A2(ext_interrupts[3]), .ZN(
        n9543) );
  NAND2_X2 U9864 ( .A1(pipeline_csr_mie[12]), .A2(ext_interrupts[4]), .ZN(
        n9542) );
  NAND2_X2 U9865 ( .A1(pipeline_csr_mie[13]), .A2(ext_interrupts[5]), .ZN(
        n9541) );
  NAND4_X2 U9866 ( .A1(n9544), .A2(n9543), .A3(n9542), .A4(n9541), .ZN(n9545)
         );
  NOR2_X2 U9867 ( .A1(n9545), .A2(n9546), .ZN(n9561) );
  NAND2_X2 U9868 ( .A1(n9547), .A2(pipeline_csr_mip_3), .ZN(n9551) );
  NAND2_X2 U9869 ( .A1(ext_interrupts[19]), .A2(n9548), .ZN(n9550) );
  NAND2_X2 U9870 ( .A1(pipeline_csr_mie[31]), .A2(ext_interrupts[23]), .ZN(
        n9549) );
  NAND3_X2 U9871 ( .A1(n9551), .A2(n9550), .A3(n9549), .ZN(n9559) );
  NAND2_X2 U9872 ( .A1(ext_interrupts[17]), .A2(n9552), .ZN(n9557) );
  NAND2_X2 U9873 ( .A1(ext_interrupts[16]), .A2(n9553), .ZN(n9556) );
  NAND2_X2 U9874 ( .A1(ext_interrupts[18]), .A2(n9554), .ZN(n9555) );
  NAND3_X2 U9875 ( .A1(n9557), .A2(n9556), .A3(n9555), .ZN(n9558) );
  NOR2_X2 U9876 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  NAND2_X2 U9877 ( .A1(ext_interrupts[9]), .A2(n9563), .ZN(n9568) );
  NAND2_X2 U9878 ( .A1(ext_interrupts[6]), .A2(n9565), .ZN(n9566) );
  NAND4_X2 U9879 ( .A1(n9569), .A2(n9567), .A3(n9568), .A4(n9566), .ZN(n9584)
         );
  NAND2_X2 U9880 ( .A1(ext_interrupts[13]), .A2(n9570), .ZN(n9574) );
  NAND2_X2 U9881 ( .A1(ext_interrupts[14]), .A2(n9571), .ZN(n9573) );
  NAND2_X2 U9882 ( .A1(ext_interrupts[12]), .A2(n10896), .ZN(n9572) );
  NAND3_X2 U9883 ( .A1(n9574), .A2(n9573), .A3(n9572), .ZN(n9583) );
  NAND2_X2 U9884 ( .A1(ext_interrupts[21]), .A2(n9575), .ZN(n9581) );
  NAND2_X2 U9885 ( .A1(ext_interrupts[22]), .A2(n9576), .ZN(n9580) );
  NAND2_X2 U9886 ( .A1(pipeline_csr_mie[7]), .A2(pipeline_csr_mip_7_), .ZN(
        n9579) );
  NAND2_X2 U9887 ( .A1(ext_interrupts[20]), .A2(n9577), .ZN(n9578) );
  NAND4_X2 U9888 ( .A1(n9581), .A2(n9580), .A3(n9579), .A4(n9578), .ZN(n9582)
         );
  NOR2_X2 U9889 ( .A1(n10323), .A2(pipeline_csr_priv_stack_0), .ZN(n9587) );
  XOR2_X2 U9890 ( .A(pipeline_ctrl_N82), .B(n10323), .Z(n9586) );
  NOR2_X2 U9891 ( .A1(ext_interrupts[6]), .A2(ext_interrupts[5]), .ZN(n9590)
         );
  NOR2_X2 U9892 ( .A1(ext_interrupts[3]), .A2(ext_interrupts[4]), .ZN(n9589)
         );
  NAND4_X2 U9893 ( .A1(n9592), .A2(n9591), .A3(n9590), .A4(n9589), .ZN(n9598)
         );
  NOR2_X2 U9894 ( .A1(ext_interrupts[19]), .A2(ext_interrupts[20]), .ZN(n9596)
         );
  NOR2_X2 U9895 ( .A1(ext_interrupts[17]), .A2(ext_interrupts[18]), .ZN(n9595)
         );
  NOR2_X2 U9896 ( .A1(ext_interrupts[14]), .A2(ext_interrupts[15]), .ZN(n9594)
         );
  NOR2_X2 U9897 ( .A1(ext_interrupts[13]), .A2(ext_interrupts[12]), .ZN(n9593)
         );
  NAND4_X2 U9898 ( .A1(n9596), .A2(n9595), .A3(n9594), .A4(n9593), .ZN(n9597)
         );
  NAND3_X2 U9899 ( .A1(n10510), .A2(n1547), .A3(n793), .ZN(n9600) );
  NOR2_X2 U9900 ( .A1(n9600), .A2(n9599), .ZN(n9604) );
  NOR2_X2 U9901 ( .A1(ext_interrupts[21]), .A2(ext_interrupts[22]), .ZN(n9603)
         );
  NOR2_X2 U9902 ( .A1(ext_interrupts[2]), .A2(ext_interrupts[1]), .ZN(n9602)
         );
  NOR2_X2 U9903 ( .A1(ext_interrupts[23]), .A2(ext_interrupts[0]), .ZN(n9601)
         );
  NAND4_X2 U9904 ( .A1(n9604), .A2(n9603), .A3(n9602), .A4(n9601), .ZN(n9606)
         );
  NOR2_X2 U9905 ( .A1(n9606), .A2(n9605), .ZN(n9612) );
  NAND2_X2 U9906 ( .A1(pipeline_md_state[1]), .A2(pipeline_md_state[0]), .ZN(
        n9608) );
  NAND2_X2 U9907 ( .A1(n9608), .A2(n9607), .ZN(n9609) );
  NAND2_X2 U9908 ( .A1(pipeline_inst_DX[0]), .A2(pipeline_inst_DX[1]), .ZN(
        n9671) );
  INV_X4 U9909 ( .A(n9671), .ZN(n12834) );
  INV_X4 U9910 ( .A(n638), .ZN(n12546) );
  NOR3_X2 U9911 ( .A1(pipeline_regfile_N16), .A2(n12546), .A3(
        pipeline_regfile_N15), .ZN(n9614) );
  NOR3_X2 U9912 ( .A1(pipeline_inst_DX[10]), .A2(pipeline_inst_DX[11]), .A3(
        n10258), .ZN(n9615) );
  NOR3_X2 U9913 ( .A1(n9650), .A2(n9631), .A3(n9651), .ZN(n9616) );
  NAND3_X2 U9914 ( .A1(n9623), .A2(n9648), .A3(n9616), .ZN(n10131) );
  INV_X4 U9915 ( .A(n10131), .ZN(n13096) );
  NAND2_X2 U9916 ( .A1(n7172), .A2(n6711), .ZN(n10237) );
  NOR3_X2 U9917 ( .A1(pipeline_inst_DX[30]), .A2(n10237), .A3(pipeline_imm_31_), .ZN(n9617) );
  NAND2_X2 U9918 ( .A1(n702), .A2(n7182), .ZN(n9619) );
  INV_X4 U9919 ( .A(n9619), .ZN(n9618) );
  NAND2_X2 U9920 ( .A1(n602), .A2(n601), .ZN(n13095) );
  INV_X4 U9921 ( .A(n13095), .ZN(n10194) );
  NAND2_X2 U9922 ( .A1(n603), .A2(n10194), .ZN(n9686) );
  INV_X4 U9923 ( .A(n9686), .ZN(n10132) );
  NAND2_X2 U9924 ( .A1(n10194), .A2(pipeline_dmem_type_2_), .ZN(n10184) );
  NAND3_X2 U9925 ( .A1(n10132), .A2(n6794), .A3(n9619), .ZN(n9620) );
  INV_X4 U9926 ( .A(n693), .ZN(n10333) );
  NOR2_X2 U9927 ( .A1(n9621), .A2(n10333), .ZN(n9622) );
  OAI22_X2 U9928 ( .A1(pipeline_inst_DX[28]), .A2(n9658), .B1(n9622), .B2(
        n9634), .ZN(n9630) );
  NAND2_X2 U9929 ( .A1(n9631), .A2(pipeline_inst_DX[2]), .ZN(n9637) );
  OAI22_X2 U9930 ( .A1(n9651), .A2(n9648), .B1(n9637), .B2(pipeline_inst_DX[3]), .ZN(n9627) );
  NOR2_X2 U9931 ( .A1(n9631), .A2(n9623), .ZN(n9624) );
  NOR2_X2 U9932 ( .A1(n9651), .A2(n9624), .ZN(n9625) );
  NOR2_X2 U9933 ( .A1(n9650), .A2(n9625), .ZN(n9626) );
  AOI221_X2 U9934 ( .B1(n9637), .B2(pipeline_inst_DX[3]), .C1(n9627), .C2(
        n9650), .A(n9626), .ZN(n9628) );
  INV_X4 U9935 ( .A(pipeline_csr_system_wen), .ZN(n4201) );
  NOR3_X2 U9936 ( .A1(n713), .A2(n10242), .A3(n4201), .ZN(n9629) );
  NAND4_X2 U9937 ( .A1(pipeline_inst_DX[6]), .A2(n9623), .A3(n9648), .A4(n7173), .ZN(n9698) );
  INV_X4 U9938 ( .A(n9698), .ZN(n12402) );
  NAND3_X2 U9939 ( .A1(pipeline_inst_DX[2]), .A2(n9648), .A3(n7173), .ZN(
        n12394) );
  NAND2_X2 U9940 ( .A1(n713), .A2(n9632), .ZN(n10246) );
  INV_X4 U9941 ( .A(n10246), .ZN(n9633) );
  NAND3_X2 U9942 ( .A1(n7086), .A2(n6794), .A3(n603), .ZN(n9636) );
  NAND2_X2 U9943 ( .A1(n7078), .A2(n702), .ZN(n13102) );
  INV_X4 U9944 ( .A(n13102), .ZN(n10248) );
  NOR2_X2 U9945 ( .A1(n7180), .A2(n601), .ZN(n9635) );
  NOR3_X2 U9946 ( .A1(n9636), .A2(dmem_hsize[1]), .A3(n9635), .ZN(n9638) );
  INV_X4 U9947 ( .A(n9637), .ZN(n9678) );
  NAND4_X2 U9948 ( .A1(n9651), .A2(pipeline_inst_DX[3]), .A3(n9678), .A4(n9650), .ZN(n9670) );
  OAI22_X2 U9949 ( .A1(n10132), .A2(n12394), .B1(n9638), .B2(n9670), .ZN(n9639) );
  AOI221_X2 U9950 ( .B1(n12402), .B2(n6795), .C1(n7083), .C2(n7075), .A(n9639), 
        .ZN(n9640) );
  NAND2_X2 U9951 ( .A1(n9641), .A2(n9640), .ZN(n11187) );
  OR3_X1 U9952 ( .A1(n7083), .A2(n11187), .A3(pipeline_ctrl_had_ex_DX), .ZN(
        n10093) );
  INV_X4 U9953 ( .A(n10093), .ZN(n10127) );
  NAND3_X2 U9954 ( .A1(pipeline_inst_DX[5]), .A2(n9623), .A3(n7080), .ZN(n9695) );
  INV_X4 U9955 ( .A(n9695), .ZN(n9643) );
  NAND2_X2 U9956 ( .A1(n7085), .A2(n12834), .ZN(n12836) );
  XNOR2_X2 U9957 ( .A(pipeline_regfile_N14), .B(pipeline_reg_to_wr_WB[2]), 
        .ZN(n9644) );
  XNOR2_X2 U9958 ( .A(n12992), .B(pipeline_regfile_N16), .ZN(n9656) );
  NAND3_X2 U9959 ( .A1(n9651), .A2(n9623), .A3(n7080), .ZN(n9704) );
  NAND2_X2 U9960 ( .A1(n9704), .A2(n9695), .ZN(n9694) );
  NAND4_X2 U9961 ( .A1(n9650), .A2(n9623), .A3(n9648), .A4(n7173), .ZN(n9666)
         );
  INV_X4 U9962 ( .A(n9666), .ZN(n10139) );
  NOR3_X2 U9963 ( .A1(pipeline_inst_DX[3]), .A2(pipeline_inst_DX[2]), .A3(
        pipeline_inst_DX[4]), .ZN(n9649) );
  NAND3_X2 U9964 ( .A1(n9651), .A2(n9650), .A3(n9649), .ZN(n10129) );
  INV_X4 U9965 ( .A(n10129), .ZN(n12835) );
  NOR2_X2 U9966 ( .A1(n10139), .A2(n12835), .ZN(n9652) );
  NAND4_X2 U9967 ( .A1(n10130), .A2(n6740), .A3(n12394), .A4(n9698), .ZN(n9655) );
  NAND3_X2 U9968 ( .A1(n10348), .A2(n6369), .A3(
        pipeline_ctrl_wr_reg_unkilled_WB), .ZN(n9667) );
  INV_X4 U9969 ( .A(n10258), .ZN(n9653) );
  NOR2_X2 U9970 ( .A1(n9667), .A2(n9653), .ZN(n9654) );
  NAND3_X2 U9971 ( .A1(n9656), .A2(n9655), .A3(n9654), .ZN(n9657) );
  XOR2_X2 U9972 ( .A(pipeline_regfile_N19), .B(n12988), .Z(n9662) );
  XOR2_X2 U9973 ( .A(n8223), .B(n12995), .Z(n9661) );
  XOR2_X2 U9974 ( .A(n693), .B(n12990), .Z(n9660) );
  XOR2_X2 U9975 ( .A(n9658), .B(pipeline_reg_to_wr_WB[1]), .Z(n9659) );
  NAND4_X2 U9976 ( .A1(n9662), .A2(n9661), .A3(n9660), .A4(n9659), .ZN(n9665)
         );
  NAND2_X2 U9977 ( .A1(n7167), .A2(n7078), .ZN(n9703) );
  INV_X4 U9978 ( .A(n9703), .ZN(n9664) );
  XOR2_X2 U9979 ( .A(pipeline_regfile_N21), .B(n12992), .Z(n9663) );
  NOR4_X2 U9980 ( .A1(n9665), .A2(n9664), .A3(n9663), .A4(n9671), .ZN(n9669)
         );
  NAND3_X2 U9981 ( .A1(n9695), .A2(n9698), .A3(n9666), .ZN(n9668) );
  NAND2_X2 U9982 ( .A1(pipeline_ctrl_dmem_en_WB), .A2(n790), .ZN(n9723) );
  NAND3_X2 U9983 ( .A1(n602), .A2(n603), .A3(dmem_hsize[0]), .ZN(n10185) );
  NOR3_X2 U9984 ( .A1(n9671), .A2(n9670), .A3(n10185), .ZN(n9672) );
  NAND3_X2 U9985 ( .A1(n7180), .A2(n9673), .A3(n9672), .ZN(n10306) );
  OAI221_X2 U9986 ( .B1(n7183), .B2(n12836), .C1(n9674), .C2(n9723), .A(n10306), .ZN(n9675) );
  NAND2_X2 U9987 ( .A1(n6743), .A2(n9675), .ZN(n9676) );
  INV_X4 U9988 ( .A(n12395), .ZN(n10092) );
  NAND2_X2 U9989 ( .A1(n10092), .A2(n13130), .ZN(n9677) );
  INV_X4 U9990 ( .A(n9677), .ZN(n12832) );
  NAND2_X2 U9991 ( .A1(n9677), .A2(n13130), .ZN(n12823) );
  INV_X4 U9992 ( .A(imem_hresp), .ZN(n10096) );
  NAND2_X2 U9993 ( .A1(n10092), .A2(n6743), .ZN(n10346) );
  INV_X4 U9994 ( .A(n10346), .ZN(n13097) );
  NAND3_X2 U9995 ( .A1(n7078), .A2(n6745), .A3(n13097), .ZN(n12396) );
  NAND3_X2 U9996 ( .A1(pipeline_inst_DX[6]), .A2(pipeline_inst_DX[5]), .A3(
        n9678), .ZN(n9722) );
  INV_X4 U9997 ( .A(n9722), .ZN(n10134) );
  NAND2_X2 U9998 ( .A1(n10134), .A2(n13097), .ZN(n9679) );
  NAND2_X2 U9999 ( .A1(n12396), .A2(n9679), .ZN(n12405) );
  INV_X4 U10000 ( .A(n12405), .ZN(n10091) );
  NAND2_X2 U10001 ( .A1(n12834), .A2(n9694), .ZN(n9691) );
  NAND2_X2 U10002 ( .A1(n12402), .A2(n12834), .ZN(n9689) );
  OAI22_X2 U10003 ( .A1(n9680), .A2(n9691), .B1(n603), .B2(n9689), .ZN(n9693)
         );
  INV_X4 U10004 ( .A(n9693), .ZN(n10082) );
  INV_X4 U10005 ( .A(n10185), .ZN(n9681) );
  NAND2_X2 U10006 ( .A1(n6738), .A2(dmem_hsize[0]), .ZN(n9688) );
  INV_X4 U10007 ( .A(n9688), .ZN(n9682) );
  NOR3_X2 U10008 ( .A1(n6784), .A2(n9681), .A3(n9682), .ZN(n9685) );
  NOR2_X2 U10009 ( .A1(dmem_hsize[1]), .A2(n601), .ZN(n9683) );
  NOR2_X2 U10010 ( .A1(n9683), .A2(n9682), .ZN(n9684) );
  OAI22_X2 U10011 ( .A1(n9685), .A2(n9691), .B1(n9684), .B2(n9689), .ZN(n9800)
         );
  NOR2_X2 U10012 ( .A1(n9686), .A2(n9695), .ZN(n9687) );
  NAND2_X2 U10013 ( .A1(n603), .A2(n601), .ZN(n9696) );
  AOI221_X2 U10014 ( .B1(n9687), .B2(pipeline_inst_DX[30]), .C1(n9696), .C2(
        dmem_hsize[1]), .A(n6741), .ZN(n9692) );
  NAND2_X2 U10015 ( .A1(n6738), .A2(n601), .ZN(n10186) );
  NAND2_X2 U10016 ( .A1(n10186), .A2(n9688), .ZN(n10193) );
  INV_X4 U10017 ( .A(n10193), .ZN(n9690) );
  OAI22_X2 U10018 ( .A1(n9692), .A2(n9691), .B1(n9690), .B2(n9689), .ZN(n10083) );
  NAND2_X2 U10019 ( .A1(n7068), .A2(n10083), .ZN(n12791) );
  INV_X4 U10020 ( .A(n10083), .ZN(n10074) );
  INV_X4 U10021 ( .A(n9694), .ZN(n10130) );
  NOR3_X2 U10022 ( .A1(n9696), .A2(n713), .A3(n9695), .ZN(n9697) );
  NOR3_X2 U10023 ( .A1(n6741), .A2(n6795), .A3(n9697), .ZN(n9699) );
  OAI22_X2 U10024 ( .A1(n10130), .A2(n9699), .B1(n6795), .B2(n9698), .ZN(n9700) );
  NAND2_X2 U10025 ( .A1(n12834), .A2(n9700), .ZN(n10085) );
  NAND3_X2 U10026 ( .A1(n6578), .A2(n9800), .A3(n10085), .ZN(n12794) );
  NAND2_X2 U10027 ( .A1(n12791), .A2(n12794), .ZN(n11159) );
  INV_X4 U10028 ( .A(n11159), .ZN(n12376) );
  NAND2_X2 U10029 ( .A1(n10139), .A2(n12834), .ZN(n9795) );
  NAND2_X2 U10030 ( .A1(n9534), .A2(pipeline_wb_src_sel_WB_0_), .ZN(n12839) );
  NAND2_X2 U10031 ( .A1(n9781), .A2(pipeline_md_resp_result[3]), .ZN(n9701) );
  OAI221_X2 U10032 ( .B1(n414), .B2(n6694), .C1(n474), .C2(n9534), .A(n9701), 
        .ZN(n9702) );
  INV_X4 U10033 ( .A(n9702), .ZN(n12967) );
  NAND2_X2 U10034 ( .A1(n7080), .A2(pipeline_inst_DX[2]), .ZN(n10128) );
  NAND3_X2 U10035 ( .A1(n6740), .A2(n9704), .A3(n10128), .ZN(n9797) );
  INV_X4 U10036 ( .A(n9797), .ZN(n10057) );
  NAND2_X2 U10037 ( .A1(n10057), .A2(n9722), .ZN(n10056) );
  INV_X4 U10038 ( .A(n10128), .ZN(n9721) );
  NAND2_X2 U10039 ( .A1(n9721), .A2(n12834), .ZN(n10044) );
  NAND2_X2 U10040 ( .A1(n9795), .A2(n9396), .ZN(n9796) );
  INV_X4 U10041 ( .A(n9796), .ZN(n9705) );
  INV_X4 U10042 ( .A(n9710), .ZN(n9790) );
  NAND2_X2 U10043 ( .A1(n9790), .A2(pipeline_regfile_N20), .ZN(n9706) );
  INV_X4 U10044 ( .A(n9795), .ZN(n9712) );
  NAND2_X2 U10045 ( .A1(n9781), .A2(pipeline_md_resp_result[2]), .ZN(n9708) );
  OAI221_X2 U10046 ( .B1(n412), .B2(n6694), .C1(n473), .C2(n9534), .A(n9708), 
        .ZN(n9709) );
  INV_X4 U10047 ( .A(n9709), .ZN(n12972) );
  OAI22_X2 U10048 ( .A1(n12972), .A2(n10055), .B1(n7096), .B2(n7061), .ZN(
        pipeline_rs2_data_bypassed[2]) );
  OAI22_X2 U10049 ( .A1(n9722), .A2(n9797), .B1(n702), .B2(n9710), .ZN(n9711)
         );
  NAND2_X2 U10050 ( .A1(n9781), .A2(pipeline_md_resp_result[1]), .ZN(n9713) );
  OAI221_X2 U10051 ( .B1(n410), .B2(n6694), .C1(n12936), .C2(n9534), .A(n9713), 
        .ZN(n9714) );
  INV_X4 U10052 ( .A(n9714), .ZN(n12977) );
  OAI22_X2 U10053 ( .A1(n12977), .A2(n6638), .B1(n7061), .B2(n7144), .ZN(
        pipeline_rs2_data_bypassed[1]) );
  INV_X4 U10054 ( .A(pipeline_rs2_data_bypassed[1]), .ZN(n9716) );
  NAND2_X2 U10055 ( .A1(n9781), .A2(pipeline_md_resp_result[0]), .ZN(n9717) );
  OAI221_X2 U10056 ( .B1(n408), .B2(n6694), .C1(n12937), .C2(n9534), .A(n9717), 
        .ZN(n9718) );
  INV_X4 U10057 ( .A(n9718), .ZN(n12987) );
  INV_X4 U10058 ( .A(pipeline_rs2_data_bypassed[0]), .ZN(n9720) );
  INV_X4 U10059 ( .A(n6617), .ZN(n11404) );
  NAND2_X2 U10060 ( .A1(n12834), .A2(n6792), .ZN(n9786) );
  NAND2_X2 U10061 ( .A1(n9781), .A2(pipeline_md_resp_result[26]), .ZN(n9725)
         );
  OAI221_X2 U10062 ( .B1(n460), .B2(n6694), .C1(n497), .C2(n9534), .A(n9725), 
        .ZN(n9726) );
  INV_X4 U10063 ( .A(n9726), .ZN(n12862) );
  OAI22_X2 U10064 ( .A1(n9440), .A2(n7116), .B1(n12862), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[26]) );
  INV_X4 U10065 ( .A(pipeline_rs1_data_bypassed[26]), .ZN(n12434) );
  NAND2_X2 U10066 ( .A1(n9786), .A2(n9397), .ZN(n9785) );
  NAND2_X2 U10067 ( .A1(n12276), .A2(n6561), .ZN(n12211) );
  NAND2_X2 U10068 ( .A1(n9781), .A2(pipeline_md_resp_result[25]), .ZN(n9727)
         );
  OAI221_X2 U10069 ( .B1(n458), .B2(n6694), .C1(n496), .C2(n9534), .A(n9727), 
        .ZN(n9728) );
  INV_X4 U10070 ( .A(n9728), .ZN(n12864) );
  OAI22_X2 U10071 ( .A1(n9439), .A2(n7105), .B1(n12864), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[25]) );
  INV_X4 U10072 ( .A(pipeline_rs1_data_bypassed[25]), .ZN(n12438) );
  NAND2_X2 U10073 ( .A1(n9471), .A2(n6609), .ZN(n12097) );
  NAND2_X2 U10074 ( .A1(n9781), .A2(pipeline_md_resp_result[24]), .ZN(n9729)
         );
  OAI221_X2 U10075 ( .B1(n456), .B2(n6694), .C1(n495), .C2(n9534), .A(n9729), 
        .ZN(n9730) );
  INV_X4 U10076 ( .A(n9730), .ZN(n12867) );
  OAI22_X2 U10077 ( .A1(n9439), .A2(n7107), .B1(n12867), .B2(n9392), .ZN(
        pipeline_rs1_data_bypassed[24]) );
  INV_X4 U10078 ( .A(pipeline_rs1_data_bypassed[24]), .ZN(n12442) );
  OAI22_X2 U10079 ( .A1(n739), .A2(n9445), .B1(n12442), .B2(n9443), .ZN(
        pipeline_alu_src_a[24]) );
  NAND2_X2 U10080 ( .A1(n9489), .A2(pipeline_alu_src_a[24]), .ZN(n11958) );
  NAND2_X2 U10081 ( .A1(n9781), .A2(pipeline_md_resp_result[27]), .ZN(n9731)
         );
  OAI221_X2 U10082 ( .B1(n462), .B2(n6694), .C1(n498), .C2(n10144), .A(n9731), 
        .ZN(n9732) );
  INV_X4 U10083 ( .A(n9732), .ZN(n12860) );
  OAI22_X2 U10084 ( .A1(n6970), .A2(n6788), .B1(n12860), .B2(n9784), .ZN(
        pipeline_rs1_data_bypassed[27]) );
  INV_X4 U10085 ( .A(pipeline_rs1_data_bypassed[27]), .ZN(n12430) );
  OAI22_X2 U10086 ( .A1(n742), .A2(n9445), .B1(n12430), .B2(n9443), .ZN(
        pipeline_alu_src_a[27]) );
  NAND4_X2 U10087 ( .A1(n12211), .A2(n12097), .A3(n11958), .A4(n12651), .ZN(
        n11952) );
  INV_X4 U10088 ( .A(n12582), .ZN(n12780) );
  NAND2_X2 U10089 ( .A1(n9781), .A2(pipeline_md_resp_result[30]), .ZN(n9733)
         );
  OAI221_X2 U10090 ( .B1(n468), .B2(n6694), .C1(n501), .C2(n9534), .A(n9733), 
        .ZN(n9734) );
  INV_X4 U10091 ( .A(n9734), .ZN(n12854) );
  OAI22_X2 U10092 ( .A1(n9440), .A2(n7115), .B1(n12854), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[30]) );
  INV_X4 U10093 ( .A(pipeline_rs1_data_bypassed[30]), .ZN(n12418) );
  NAND2_X2 U10094 ( .A1(n12276), .A2(n6997), .ZN(n9742) );
  NAND2_X2 U10095 ( .A1(n9781), .A2(pipeline_md_resp_result[29]), .ZN(n9735)
         );
  OAI221_X2 U10096 ( .B1(n466), .B2(n6694), .C1(n500), .C2(n9534), .A(n9735), 
        .ZN(n9736) );
  INV_X4 U10097 ( .A(n9736), .ZN(n12856) );
  OAI22_X2 U10098 ( .A1(n9439), .A2(n7114), .B1(n12856), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[29]) );
  INV_X4 U10099 ( .A(pipeline_rs1_data_bypassed[29]), .ZN(n12422) );
  NAND2_X2 U10100 ( .A1(n9471), .A2(pipeline_alu_src_a[29]), .ZN(n12653) );
  NAND2_X2 U10101 ( .A1(n9781), .A2(pipeline_md_resp_result[28]), .ZN(n9737)
         );
  OAI221_X2 U10102 ( .B1(n464), .B2(n6694), .C1(n499), .C2(n10144), .A(n9737), 
        .ZN(n9738) );
  INV_X4 U10103 ( .A(n9738), .ZN(n12858) );
  OAI22_X2 U10104 ( .A1(n9440), .A2(n7117), .B1(n12858), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[28]) );
  INV_X4 U10105 ( .A(pipeline_rs1_data_bypassed[28]), .ZN(n12426) );
  NAND2_X2 U10106 ( .A1(n9489), .A2(n6565), .ZN(n12209) );
  NAND2_X2 U10107 ( .A1(n9781), .A2(pipeline_md_resp_result[31]), .ZN(n9739)
         );
  OAI221_X2 U10108 ( .B1(n470), .B2(n6694), .C1(n502), .C2(n9534), .A(n9739), 
        .ZN(n9740) );
  INV_X4 U10109 ( .A(n9740), .ZN(n12852) );
  OAI22_X2 U10110 ( .A1(n9439), .A2(n7101), .B1(n12852), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[31]) );
  NAND2_X2 U10111 ( .A1(n11869), .A2(n7006), .ZN(n9741) );
  NAND4_X2 U10112 ( .A1(n9742), .A2(n12653), .A3(n12209), .A4(n9741), .ZN(
        n12208) );
  NAND2_X2 U10113 ( .A1(n9781), .A2(pipeline_md_resp_result[18]), .ZN(n9743)
         );
  OAI221_X2 U10114 ( .B1(n444), .B2(n6694), .C1(n489), .C2(n10144), .A(n9743), 
        .ZN(n12885) );
  INV_X4 U10115 ( .A(n12885), .ZN(n9954) );
  INV_X4 U10116 ( .A(pipeline_rs1_data_bypassed[18]), .ZN(n12466) );
  NAND2_X2 U10117 ( .A1(n12276), .A2(pipeline_alu_src_a[18]), .ZN(n11619) );
  NAND2_X2 U10118 ( .A1(n9781), .A2(pipeline_md_resp_result[17]), .ZN(n9744)
         );
  OAI221_X2 U10119 ( .B1(n442), .B2(n6694), .C1(n488), .C2(n10144), .A(n9744), 
        .ZN(n12888) );
  INV_X4 U10120 ( .A(n12888), .ZN(n9819) );
  NAND2_X2 U10121 ( .A1(n9781), .A2(pipeline_md_resp_result[16]), .ZN(n9745)
         );
  OAI221_X2 U10122 ( .B1(n440), .B2(n6694), .C1(n487), .C2(n10144), .A(n9745), 
        .ZN(n12894) );
  INV_X4 U10123 ( .A(n12894), .ZN(n9825) );
  INV_X4 U10124 ( .A(pipeline_rs1_data_bypassed[16]), .ZN(n12474) );
  OAI22_X2 U10125 ( .A1(n731), .A2(n9445), .B1(n12474), .B2(n9443), .ZN(
        pipeline_alu_src_a[16]) );
  NAND2_X2 U10126 ( .A1(n9781), .A2(pipeline_md_resp_result[19]), .ZN(n9746)
         );
  OAI221_X2 U10127 ( .B1(n446), .B2(n6694), .C1(n490), .C2(n10144), .A(n9746), 
        .ZN(n12882) );
  INV_X4 U10128 ( .A(n12882), .ZN(n9966) );
  OAI22_X2 U10129 ( .A1(n9440), .A2(n7113), .B1(n9966), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[19]) );
  INV_X4 U10130 ( .A(pipeline_rs1_data_bypassed[19]), .ZN(n12462) );
  NAND2_X2 U10131 ( .A1(n11869), .A2(pipeline_alu_src_a[19]), .ZN(n11774) );
  NAND4_X2 U10132 ( .A1(n11619), .A2(n9748), .A3(n9747), .A4(n11774), .ZN(
        n12779) );
  INV_X4 U10133 ( .A(n12779), .ZN(n11643) );
  NAND2_X2 U10134 ( .A1(n9781), .A2(pipeline_md_resp_result[22]), .ZN(n9749)
         );
  OAI221_X2 U10135 ( .B1(n452), .B2(n6694), .C1(n493), .C2(n10144), .A(n9749), 
        .ZN(n12873) );
  INV_X4 U10136 ( .A(n12873), .ZN(n9985) );
  INV_X4 U10137 ( .A(pipeline_rs1_data_bypassed[22]), .ZN(n12450) );
  OAI22_X2 U10138 ( .A1(n737), .A2(n9445), .B1(n12450), .B2(n9443), .ZN(
        pipeline_alu_src_a[22]) );
  NAND2_X2 U10139 ( .A1(n12276), .A2(n6626), .ZN(n11960) );
  NAND2_X2 U10140 ( .A1(n9781), .A2(pipeline_md_resp_result[21]), .ZN(n9750)
         );
  OAI221_X2 U10141 ( .B1(n450), .B2(n6694), .C1(n492), .C2(n10144), .A(n9750), 
        .ZN(n12876) );
  INV_X4 U10142 ( .A(n12876), .ZN(n9814) );
  OAI22_X2 U10143 ( .A1(n9439), .A2(n7110), .B1(n9814), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[21]) );
  INV_X4 U10144 ( .A(pipeline_rs1_data_bypassed[21]), .ZN(n12454) );
  OAI22_X2 U10145 ( .A1(n736), .A2(n9445), .B1(n12454), .B2(n9443), .ZN(
        pipeline_alu_src_a[21]) );
  NAND2_X2 U10146 ( .A1(n9471), .A2(pipeline_alu_src_a[21]), .ZN(n11776) );
  NAND2_X2 U10147 ( .A1(n9781), .A2(pipeline_md_resp_result[20]), .ZN(n9751)
         );
  OAI221_X2 U10148 ( .B1(n448), .B2(n6694), .C1(n491), .C2(n10144), .A(n9751), 
        .ZN(n12879) );
  INV_X4 U10149 ( .A(n12879), .ZN(n9811) );
  OAI22_X2 U10150 ( .A1(n9439), .A2(n7111), .B1(n9811), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[20]) );
  INV_X4 U10151 ( .A(pipeline_rs1_data_bypassed[20]), .ZN(n12458) );
  OAI22_X2 U10152 ( .A1(n735), .A2(n9445), .B1(n12458), .B2(n9443), .ZN(
        pipeline_alu_src_a[20]) );
  NAND2_X2 U10153 ( .A1(n9489), .A2(pipeline_alu_src_a[20]), .ZN(n11617) );
  NAND2_X2 U10154 ( .A1(n9781), .A2(pipeline_md_resp_result[23]), .ZN(n9752)
         );
  INV_X4 U10156 ( .A(n12870), .ZN(n9997) );
  OAI22_X2 U10157 ( .A1(n9440), .A2(n7109), .B1(n9997), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[23]) );
  OAI22_X2 U10158 ( .A1(n738), .A2(n9445), .B1(n12446), .B2(n9443), .ZN(
        pipeline_alu_src_a[23]) );
  NAND2_X2 U10159 ( .A1(n11869), .A2(n6980), .ZN(n12095) );
  NAND4_X2 U10160 ( .A1(n11960), .A2(n11776), .A3(n11617), .A4(n12095), .ZN(
        n11985) );
  INV_X4 U10161 ( .A(n11985), .ZN(n11607) );
  OAI22_X2 U10162 ( .A1(n11643), .A2(n9509), .B1(n11607), .B2(n12774), .ZN(
        n9753) );
  AOI221_X2 U10163 ( .B1(n9511), .B2(n11952), .C1(n12780), .C2(n12208), .A(
        n9753), .ZN(n11378) );
  NAND2_X2 U10164 ( .A1(n9781), .A2(pipeline_md_resp_result[9]), .ZN(n9754) );
  INV_X4 U10166 ( .A(n9755), .ZN(n12933) );
  NAND2_X2 U10167 ( .A1(n9781), .A2(pipeline_md_resp_result[10]), .ZN(n9756)
         );
  OAI221_X2 U10168 ( .B1(n428), .B2(n6694), .C1(n481), .C2(n10144), .A(n9756), 
        .ZN(n9757) );
  INV_X4 U10169 ( .A(n9757), .ZN(n12928) );
  OAI22_X2 U10170 ( .A1(n9440), .A2(n7121), .B1(n12928), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[10]) );
  INV_X4 U10171 ( .A(pipeline_rs1_data_bypassed[10]), .ZN(n12497) );
  NAND2_X2 U10172 ( .A1(n9781), .A2(pipeline_md_resp_result[8]), .ZN(n9758) );
  OAI221_X2 U10173 ( .B1(n424), .B2(n6694), .C1(n479), .C2(n10144), .A(n9758), 
        .ZN(n9759) );
  INV_X4 U10174 ( .A(n9759), .ZN(n12941) );
  OAI22_X2 U10175 ( .A1(n9439), .A2(n7140), .B1(n9393), .B2(n12941), .ZN(
        pipeline_rs1_data_bypassed[8]) );
  INV_X4 U10176 ( .A(pipeline_rs1_data_bypassed[8]), .ZN(n12505) );
  NAND2_X2 U10177 ( .A1(n9781), .A2(pipeline_md_resp_result[11]), .ZN(n9760)
         );
  OAI221_X2 U10178 ( .B1(n430), .B2(n6694), .C1(n482), .C2(n10144), .A(n9760), 
        .ZN(n9761) );
  INV_X4 U10179 ( .A(n9761), .ZN(n12923) );
  OAI22_X2 U10180 ( .A1(n9440), .A2(n7146), .B1(n12923), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[11]) );
  INV_X4 U10181 ( .A(pipeline_rs1_data_bypassed[11]), .ZN(n12493) );
  OAI22_X2 U10182 ( .A1(n9334), .A2(n12565), .B1(n6613), .B2(n9401), .ZN(n9762) );
  NAND2_X2 U10183 ( .A1(n9781), .A2(pipeline_md_resp_result[13]), .ZN(n9763)
         );
  OAI221_X2 U10184 ( .B1(n434), .B2(n6694), .C1(n484), .C2(n10144), .A(n9763), 
        .ZN(n9764) );
  INV_X4 U10185 ( .A(n9764), .ZN(n12913) );
  OAI22_X2 U10186 ( .A1(n9440), .A2(n7103), .B1(n12913), .B2(n9784), .ZN(
        pipeline_rs1_data_bypassed[13]) );
  INV_X4 U10187 ( .A(pipeline_rs1_data_bypassed[13]), .ZN(n12485) );
  OAI22_X2 U10188 ( .A1(n728), .A2(n9445), .B1(n12485), .B2(n9443), .ZN(
        pipeline_alu_src_a[13]) );
  NAND2_X2 U10189 ( .A1(n9781), .A2(pipeline_md_resp_result[14]), .ZN(n9765)
         );
  OAI221_X2 U10190 ( .B1(n436), .B2(n6694), .C1(n485), .C2(n10144), .A(n9765), 
        .ZN(n9766) );
  INV_X4 U10191 ( .A(n9766), .ZN(n12908) );
  OAI22_X2 U10192 ( .A1(n6970), .A2(n7092), .B1(n12908), .B2(n9441), .ZN(
        pipeline_rs1_data_bypassed[14]) );
  INV_X4 U10193 ( .A(pipeline_rs1_data_bypassed[14]), .ZN(n12481) );
  NAND2_X2 U10194 ( .A1(n9781), .A2(pipeline_md_resp_result[12]), .ZN(n9767)
         );
  OAI221_X2 U10195 ( .B1(n432), .B2(n6694), .C1(n483), .C2(n10144), .A(n9767), 
        .ZN(n9768) );
  INV_X4 U10196 ( .A(n9768), .ZN(n12918) );
  OAI22_X2 U10197 ( .A1(n9439), .A2(n7142), .B1(n12918), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[12]) );
  INV_X4 U10198 ( .A(pipeline_rs1_data_bypassed[12]), .ZN(n12489) );
  NAND2_X2 U10199 ( .A1(n9781), .A2(pipeline_md_resp_result[15]), .ZN(n9769)
         );
  OAI221_X2 U10200 ( .B1(n438), .B2(n6694), .C1(n486), .C2(n10144), .A(n9769), 
        .ZN(n9770) );
  INV_X4 U10201 ( .A(n9770), .ZN(n12904) );
  OAI22_X2 U10202 ( .A1(n9440), .A2(n7099), .B1(n12904), .B2(n9393), .ZN(
        pipeline_rs1_data_bypassed[15]) );
  INV_X4 U10203 ( .A(pipeline_rs1_data_bypassed[15]), .ZN(n12477) );
  AOI221_X2 U10204 ( .B1(n9471), .B2(n6567), .C1(n12276), .C2(
        pipeline_alu_src_a[14]), .A(n9771), .ZN(n12773) );
  OAI22_X2 U10205 ( .A1(n9338), .A2(n7138), .B1(n12972), .B2(n9784), .ZN(
        pipeline_rs1_data_bypassed[2]) );
  INV_X4 U10206 ( .A(pipeline_rs1_data_bypassed[2]), .ZN(n12530) );
  NAND2_X2 U10207 ( .A1(n9471), .A2(n6632), .ZN(n9772) );
  NAND2_X2 U10208 ( .A1(n9510), .A2(n9773), .ZN(n9774) );
  OAI221_X2 U10209 ( .B1(n12775), .B2(n12645), .C1(n12773), .C2(n12582), .A(
        n9774), .ZN(n9789) );
  NAND2_X2 U10210 ( .A1(n9781), .A2(pipeline_md_resp_result[5]), .ZN(n9775) );
  OAI221_X2 U10211 ( .B1(n418), .B2(n6694), .C1(n476), .C2(n10144), .A(n9775), 
        .ZN(n9776) );
  INV_X4 U10212 ( .A(n9776), .ZN(n12957) );
  NAND2_X2 U10213 ( .A1(n9781), .A2(pipeline_md_resp_result[6]), .ZN(n9777) );
  OAI221_X2 U10214 ( .B1(n420), .B2(n6694), .C1(n477), .C2(n10144), .A(n9777), 
        .ZN(n9778) );
  INV_X4 U10215 ( .A(n9778), .ZN(n12952) );
  OAI22_X2 U10216 ( .A1(n9440), .A2(n7141), .B1(n12952), .B2(n9392), .ZN(
        pipeline_rs1_data_bypassed[6]) );
  INV_X4 U10217 ( .A(pipeline_rs1_data_bypassed[6]), .ZN(n12513) );
  NAND2_X2 U10218 ( .A1(n9781), .A2(pipeline_md_resp_result[4]), .ZN(n9779) );
  INV_X4 U10220 ( .A(n9780), .ZN(n12962) );
  NAND2_X2 U10221 ( .A1(n9781), .A2(pipeline_md_resp_result[7]), .ZN(n9782) );
  INV_X4 U10223 ( .A(n12944), .ZN(n9846) );
  INV_X4 U10224 ( .A(pipeline_rs1_data_bypassed[7]), .ZN(n12509) );
  NOR2_X2 U10225 ( .A1(n12777), .A2(n9507), .ZN(n9788) );
  OAI22_X2 U10226 ( .A1(n12987), .A2(n9393), .B1(n9440), .B2(n7093), .ZN(
        pipeline_rs1_data_bypassed[0]) );
  INV_X4 U10227 ( .A(pipeline_rs1_data_bypassed[0]), .ZN(n11279) );
  INV_X4 U10228 ( .A(n11372), .ZN(n9787) );
  NOR3_X2 U10229 ( .A1(n9789), .A2(n9788), .A3(n9787), .ZN(n9793) );
  NAND2_X2 U10230 ( .A1(n9790), .A2(pipeline_regfile_N21), .ZN(n9791) );
  MUX2_X2 U10231 ( .A(n11378), .B(n9793), .S(n12800), .Z(n9794) );
  NOR2_X2 U10232 ( .A1(n12376), .A2(n9794), .ZN(n10080) );
  INV_X4 U10233 ( .A(n6565), .ZN(n12200) );
  INV_X4 U10234 ( .A(n10085), .ZN(n9801) );
  INV_X4 U10235 ( .A(n9800), .ZN(n10081) );
  OAI22_X2 U10236 ( .A1(n9447), .A2(n7136), .B1(n12858), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[28]) );
  INV_X4 U10237 ( .A(pipeline_rs2_data_bypassed[28]), .ZN(n9799) );
  NAND2_X2 U10238 ( .A1(n9796), .A2(n9795), .ZN(n9798) );
  INV_X4 U10239 ( .A(n9915), .ZN(n9820) );
  OAI221_X2 U10240 ( .B1(n9799), .B2(n9448), .C1(n9634), .C2(n10044), .A(
        n10043), .ZN(pipeline_alu_src_b[28]) );
  INV_X4 U10241 ( .A(pipeline_alu_src_b[28]), .ZN(n12202) );
  OAI22_X2 U10242 ( .A1(n12200), .A2(n9453), .B1(n12202), .B2(n9451), .ZN(
        n10035) );
  OAI22_X2 U10243 ( .A1(n12202), .A2(n9453), .B1(n12200), .B2(n9450), .ZN(
        n10037) );
  INV_X4 U10244 ( .A(n10037), .ZN(n9804) );
  INV_X4 U10245 ( .A(pipeline_alu_src_a[29]), .ZN(n12297) );
  OAI22_X2 U10246 ( .A1(n12856), .A2(n10055), .B1(n7061), .B2(n7135), .ZN(
        pipeline_rs2_data_bypassed[29]) );
  INV_X4 U10247 ( .A(pipeline_rs2_data_bypassed[29]), .ZN(n9802) );
  OAI22_X2 U10248 ( .A1(n12297), .A2(n9453), .B1(n12299), .B2(n9451), .ZN(
        n10047) );
  OAI22_X2 U10249 ( .A1(n12299), .A2(n9456), .B1(n12297), .B2(n9451), .ZN(
        n10049) );
  INV_X4 U10250 ( .A(n10049), .ZN(n9803) );
  INV_X4 U10251 ( .A(pipeline_alu_src_a[24]), .ZN(n11962) );
  OAI22_X2 U10252 ( .A1(n9447), .A2(n7127), .B1(n12867), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[24]) );
  INV_X4 U10253 ( .A(pipeline_rs2_data_bypassed[24]), .ZN(n9805) );
  INV_X4 U10254 ( .A(pipeline_alu_src_b[24]), .ZN(n9806) );
  OAI22_X2 U10255 ( .A1(n11962), .A2(n9456), .B1(n9806), .B2(n9450), .ZN(
        n10007) );
  OAI22_X2 U10256 ( .A1(n9806), .A2(n9456), .B1(n11962), .B2(n9450), .ZN(
        n10009) );
  OAI22_X2 U10257 ( .A1(n9447), .A2(n7124), .B1(n12864), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[25]) );
  INV_X4 U10258 ( .A(pipeline_rs2_data_bypassed[25]), .ZN(n9807) );
  OAI221_X2 U10259 ( .B1(n9807), .B2(n9448), .C1(n10336), .C2(n10044), .A(
        n10043), .ZN(pipeline_alu_src_b[25]) );
  INV_X4 U10260 ( .A(pipeline_alu_src_b[25]), .ZN(n9808) );
  OAI22_X2 U10261 ( .A1(n6607), .A2(n9456), .B1(n9808), .B2(n9450), .ZN(n10018) );
  OAI22_X2 U10262 ( .A1(n9808), .A2(n9456), .B1(n6607), .B2(n9450), .ZN(n10020) );
  INV_X4 U10263 ( .A(n10020), .ZN(n9809) );
  OAI22_X2 U10264 ( .A1(n7061), .A2(n7128), .B1(n9811), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[20]) );
  INV_X4 U10265 ( .A(pipeline_rs2_data_bypassed[20]), .ZN(n9812) );
  OAI221_X2 U10266 ( .B1(n9812), .B2(n9448), .C1(n693), .C2(n9396), .A(n10043), 
        .ZN(pipeline_alu_src_b[20]) );
  INV_X4 U10267 ( .A(pipeline_alu_src_b[20]), .ZN(n9813) );
  OAI22_X2 U10268 ( .A1(n6925), .A2(n9456), .B1(n9813), .B2(n9450), .ZN(n9977)
         );
  OAI22_X2 U10269 ( .A1(n9813), .A2(n9456), .B1(n6925), .B2(n9450), .ZN(n9979)
         );
  INV_X4 U10270 ( .A(n9979), .ZN(n9818) );
  INV_X4 U10271 ( .A(pipeline_alu_src_a[21]), .ZN(n11693) );
  OAI22_X2 U10272 ( .A1(n9447), .A2(n7129), .B1(n9814), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[21]) );
  INV_X4 U10273 ( .A(pipeline_rs2_data_bypassed[21]), .ZN(n9815) );
  OAI221_X2 U10274 ( .B1(n9815), .B2(n9448), .C1(n6628), .C2(n9397), .A(n10043), .ZN(pipeline_alu_src_b[21]) );
  OAI22_X2 U10275 ( .A1(n11693), .A2(n9456), .B1(n9816), .B2(n9450), .ZN(n9989) );
  OAI22_X2 U10276 ( .A1(n9816), .A2(n9456), .B1(n11693), .B2(n9450), .ZN(n9991) );
  INV_X4 U10277 ( .A(pipeline_rs2_data_bypassed[17]), .ZN(n9821) );
  OAI221_X2 U10278 ( .B1(n9821), .B2(n9448), .C1(n638), .C2(n10044), .A(n9967), 
        .ZN(pipeline_alu_src_b[17]) );
  INV_X4 U10279 ( .A(pipeline_alu_src_b[17]), .ZN(n9822) );
  OAI22_X2 U10280 ( .A1(n11546), .A2(n9456), .B1(n9822), .B2(n9450), .ZN(n9958) );
  OAI22_X2 U10281 ( .A1(n9822), .A2(n9456), .B1(n11546), .B2(n9450), .ZN(n9959) );
  NOR2_X2 U10282 ( .A1(n9960), .A2(n9959), .ZN(n9843) );
  INV_X4 U10283 ( .A(pipeline_rs2_data_bypassed[15]), .ZN(n9823) );
  OAI221_X2 U10284 ( .B1(n9823), .B2(n9448), .C1(n636), .C2(n9396), .A(n9967), 
        .ZN(pipeline_alu_src_b[15]) );
  INV_X4 U10285 ( .A(pipeline_alu_src_b[15]), .ZN(n11347) );
  OAI22_X2 U10286 ( .A1(n11414), .A2(n9456), .B1(n11347), .B2(n9450), .ZN(
        n9832) );
  INV_X4 U10287 ( .A(n9832), .ZN(n9824) );
  OAI22_X2 U10288 ( .A1(n11347), .A2(n9455), .B1(n11414), .B2(n9451), .ZN(
        n9829) );
  NAND2_X2 U10289 ( .A1(n9824), .A2(n9829), .ZN(n9948) );
  OAI22_X2 U10290 ( .A1(n7061), .A2(n7131), .B1(n9825), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[16]) );
  INV_X4 U10291 ( .A(pipeline_rs2_data_bypassed[16]), .ZN(n9826) );
  OAI221_X2 U10292 ( .B1(n9826), .B2(n9448), .C1(n637), .C2(n9397), .A(n9967), 
        .ZN(pipeline_alu_src_b[16]) );
  INV_X4 U10293 ( .A(pipeline_alu_src_b[16]), .ZN(n9827) );
  OAI22_X2 U10294 ( .A1(n11474), .A2(n9455), .B1(n9827), .B2(n9450), .ZN(n9837) );
  INV_X4 U10295 ( .A(n9837), .ZN(n9828) );
  OAI22_X2 U10296 ( .A1(n9827), .A2(n9455), .B1(n11474), .B2(n9451), .ZN(n9836) );
  NAND2_X2 U10297 ( .A1(n9828), .A2(n9836), .ZN(n9947) );
  NAND2_X2 U10298 ( .A1(n9948), .A2(n9947), .ZN(n9834) );
  INV_X4 U10299 ( .A(n9829), .ZN(n9830) );
  NAND3_X2 U10300 ( .A1(n9832), .A2(n9831), .A3(n9830), .ZN(n9841) );
  OAI22_X2 U10301 ( .A1(n7061), .A2(n7095), .B1(n12908), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[14]) );
  INV_X4 U10302 ( .A(pipeline_rs2_data_bypassed[14]), .ZN(n9833) );
  INV_X4 U10303 ( .A(pipeline_alu_src_b[14]), .ZN(n11174) );
  INV_X4 U10304 ( .A(pipeline_alu_src_a[14]), .ZN(n11570) );
  OAI22_X2 U10305 ( .A1(n11174), .A2(n9455), .B1(n11570), .B2(n9450), .ZN(
        n9944) );
  INV_X4 U10306 ( .A(n9944), .ZN(n9835) );
  OAI22_X2 U10307 ( .A1(n11570), .A2(n9455), .B1(n11174), .B2(n9451), .ZN(
        n9942) );
  NAND3_X2 U10308 ( .A1(n9835), .A2(n9831), .A3(n9942), .ZN(n9840) );
  NAND2_X2 U10309 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  NAND3_X2 U10310 ( .A1(n9841), .A2(n9840), .A3(n9839), .ZN(n9842) );
  NOR2_X2 U10311 ( .A1(n9843), .A2(n9842), .ZN(n9965) );
  OAI22_X2 U10312 ( .A1(n7061), .A2(n7098), .B1(n12952), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[6]) );
  INV_X4 U10313 ( .A(pipeline_rs2_data_bypassed[6]), .ZN(n9844) );
  OAI22_X2 U10314 ( .A1(n9844), .A2(n9448), .B1(n10338), .B2(n9915), .ZN(
        pipeline_alu_src_b[6]) );
  INV_X4 U10315 ( .A(pipeline_alu_src_b[6]), .ZN(n11809) );
  OAI22_X2 U10316 ( .A1(n6604), .A2(n9455), .B1(n11809), .B2(n9451), .ZN(n9901) );
  NAND2_X2 U10317 ( .A1(n9901), .A2(n9845), .ZN(n9854) );
  INV_X4 U10318 ( .A(pipeline_rs2_data_bypassed[7]), .ZN(n9847) );
  OAI22_X2 U10319 ( .A1(n11885), .A2(n9455), .B1(n6610), .B2(n9451), .ZN(n9850) );
  INV_X4 U10320 ( .A(n9850), .ZN(n9848) );
  OAI22_X2 U10321 ( .A1(n6610), .A2(n9455), .B1(n11885), .B2(n9450), .ZN(n9849) );
  NAND2_X2 U10322 ( .A1(n9851), .A2(n9850), .ZN(n9902) );
  INV_X4 U10323 ( .A(n9902), .ZN(n9852) );
  INV_X4 U10324 ( .A(pipeline_rs2_data_bypassed[8]), .ZN(n9855) );
  OAI22_X2 U10325 ( .A1(n9334), .A2(n9455), .B1(n9387), .B2(n9451), .ZN(n9857)
         );
  NAND2_X2 U10326 ( .A1(n9856), .A2(n9858), .ZN(n9900) );
  INV_X4 U10327 ( .A(pipeline_rs2_data_bypassed[9]), .ZN(n9859) );
  INV_X4 U10328 ( .A(pipeline_alu_src_b[9]), .ZN(n12067) );
  INV_X4 U10329 ( .A(n6972), .ZN(n12064) );
  OAI22_X2 U10330 ( .A1(n12067), .A2(n9455), .B1(n12064), .B2(n9451), .ZN(
        n9914) );
  OAI22_X2 U10331 ( .A1(n12064), .A2(n9454), .B1(n12067), .B2(n9450), .ZN(
        n9913) );
  INV_X4 U10332 ( .A(n9913), .ZN(n9860) );
  NOR2_X2 U10333 ( .A1(n9914), .A2(n9860), .ZN(n9861) );
  NOR2_X2 U10334 ( .A1(n6943), .A2(n9451), .ZN(n9866) );
  NOR2_X2 U10335 ( .A1(n6616), .A2(n9451), .ZN(n9865) );
  NOR2_X2 U10336 ( .A1(n11404), .A2(n9456), .ZN(n9864) );
  NOR3_X2 U10337 ( .A1(n9866), .A2(n9865), .A3(n9864), .ZN(n9868) );
  OAI22_X2 U10338 ( .A1(n6631), .A2(n9454), .B1(n11405), .B2(n9451), .ZN(n9869) );
  OAI22_X2 U10339 ( .A1(n11405), .A2(n9454), .B1(n6631), .B2(n9451), .ZN(n9871) );
  NAND2_X2 U10340 ( .A1(n9871), .A2(n9870), .ZN(n9878) );
  OAI22_X2 U10341 ( .A1(n12265), .A2(n9454), .B1(n12274), .B2(n9451), .ZN(
        n9881) );
  OAI22_X2 U10342 ( .A1(n12274), .A2(n9454), .B1(n12265), .B2(n9451), .ZN(
        n9884) );
  NAND2_X2 U10343 ( .A1(n9881), .A2(n9872), .ZN(n9877) );
  OAI22_X2 U10344 ( .A1(n7009), .A2(n9454), .B1(n6633), .B2(n9450), .ZN(n9888)
         );
  INV_X4 U10345 ( .A(n9883), .ZN(n9874) );
  NAND3_X2 U10346 ( .A1(n9878), .A2(n9877), .A3(n9876), .ZN(n9879) );
  NOR2_X2 U10347 ( .A1(n9880), .A2(n9879), .ZN(n9909) );
  INV_X4 U10348 ( .A(n9881), .ZN(n9886) );
  NAND2_X2 U10349 ( .A1(n9882), .A2(n9883), .ZN(n9887) );
  OAI22_X2 U10350 ( .A1(n9447), .A2(n7119), .B1(n12957), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[5]) );
  INV_X4 U10351 ( .A(pipeline_rs2_data_bypassed[5]), .ZN(n9893) );
  OAI22_X2 U10352 ( .A1(n9893), .A2(n9448), .B1(n10336), .B2(n9915), .ZN(
        pipeline_alu_src_b[5]) );
  INV_X4 U10353 ( .A(pipeline_alu_src_b[5]), .ZN(n11732) );
  OAI22_X2 U10354 ( .A1(n11732), .A2(n9454), .B1(n6619), .B2(n9451), .ZN(n9894) );
  INV_X4 U10355 ( .A(n9894), .ZN(n9904) );
  OAI22_X2 U10356 ( .A1(n6619), .A2(n9454), .B1(n11732), .B2(n9451), .ZN(n9903) );
  NOR2_X2 U10357 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  OAI22_X2 U10358 ( .A1(n7061), .A2(n7102), .B1(n12923), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[11]) );
  NAND2_X2 U10359 ( .A1(n9449), .A2(pipeline_rs2_data_bypassed[11]), .ZN(n9910) );
  NAND2_X2 U10360 ( .A1(n9967), .A2(n9910), .ZN(pipeline_alu_src_b[11]) );
  INV_X4 U10361 ( .A(pipeline_alu_src_b[11]), .ZN(n11589) );
  OAI22_X2 U10362 ( .A1(n6613), .A2(n9453), .B1(n11589), .B2(n9450), .ZN(n9927) );
  INV_X4 U10363 ( .A(n9927), .ZN(n9911) );
  OAI22_X2 U10364 ( .A1(n11589), .A2(n9453), .B1(n6613), .B2(n9450), .ZN(n9926) );
  NAND2_X2 U10365 ( .A1(n9911), .A2(n9926), .ZN(n9930) );
  INV_X4 U10366 ( .A(pipeline_rs2_data_bypassed[12]), .ZN(n9912) );
  NAND2_X2 U10367 ( .A1(n6926), .A2(n9933), .ZN(n9929) );
  OAI22_X2 U10368 ( .A1(n9447), .A2(n7094), .B1(n12928), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[10]) );
  INV_X4 U10369 ( .A(pipeline_rs2_data_bypassed[10]), .ZN(n9916) );
  INV_X4 U10370 ( .A(pipeline_alu_src_b[10]), .ZN(n11513) );
  OAI22_X2 U10371 ( .A1(n11513), .A2(n9453), .B1(n11510), .B2(n9450), .ZN(
        n9923) );
  OAI22_X2 U10372 ( .A1(n11510), .A2(n9453), .B1(n11513), .B2(n9450), .ZN(
        n9925) );
  NAND2_X2 U10373 ( .A1(n9923), .A2(n9917), .ZN(n9918) );
  NAND2_X2 U10374 ( .A1(n9919), .A2(n9918), .ZN(n9920) );
  AOI211_X4 U10375 ( .C1(n9922), .C2(n9921), .A(n9938), .B(n9920), .ZN(n9953)
         );
  INV_X4 U10376 ( .A(n9923), .ZN(n9924) );
  INV_X4 U10377 ( .A(n9926), .ZN(n9928) );
  INV_X4 U10378 ( .A(n6568), .ZN(n11573) );
  OAI22_X2 U10379 ( .A1(n9447), .A2(n7118), .B1(n12913), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[13]) );
  INV_X4 U10380 ( .A(pipeline_rs2_data_bypassed[13]), .ZN(n9931) );
  INV_X4 U10381 ( .A(pipeline_alu_src_b[13]), .ZN(n11446) );
  OAI22_X2 U10382 ( .A1(n11573), .A2(n9453), .B1(n11446), .B2(n9451), .ZN(
        n9939) );
  OAI22_X2 U10383 ( .A1(n11446), .A2(n9453), .B1(n11573), .B2(n6744), .ZN(
        n9941) );
  INV_X4 U10384 ( .A(n9941), .ZN(n9932) );
  NAND2_X2 U10385 ( .A1(n9939), .A2(n9932), .ZN(n9937) );
  NAND2_X2 U10386 ( .A1(n9935), .A2(n9934), .ZN(n9936) );
  INV_X4 U10387 ( .A(n9939), .ZN(n9940) );
  NAND2_X2 U10388 ( .A1(n9941), .A2(n9940), .ZN(n9946) );
  INV_X4 U10389 ( .A(n9942), .ZN(n9943) );
  NAND2_X2 U10390 ( .A1(n9944), .A2(n9943), .ZN(n9945) );
  NAND2_X2 U10391 ( .A1(n9946), .A2(n9945), .ZN(n9950) );
  NAND2_X2 U10392 ( .A1(n9948), .A2(n9947), .ZN(n9949) );
  NOR2_X2 U10393 ( .A1(n9950), .A2(n9949), .ZN(n9951) );
  OAI21_X4 U10394 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9964) );
  OAI22_X2 U10395 ( .A1(n7061), .A2(n7132), .B1(n9954), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[18]) );
  INV_X4 U10396 ( .A(pipeline_rs2_data_bypassed[18]), .ZN(n9955) );
  OAI221_X2 U10397 ( .B1(n9955), .B2(n10056), .C1(n9279), .C2(n10044), .A(
        n9967), .ZN(pipeline_alu_src_b[18]) );
  INV_X4 U10398 ( .A(pipeline_alu_src_b[18]), .ZN(n9956) );
  INV_X4 U10399 ( .A(pipeline_alu_src_a[18]), .ZN(n11547) );
  OAI22_X2 U10400 ( .A1(n9956), .A2(n9453), .B1(n11547), .B2(n6744), .ZN(n9971) );
  OAI22_X2 U10401 ( .A1(n11547), .A2(n9453), .B1(n9956), .B2(n6744), .ZN(n9973) );
  INV_X4 U10402 ( .A(n9973), .ZN(n9957) );
  NAND2_X2 U10403 ( .A1(n9971), .A2(n9957), .ZN(n9962) );
  INV_X4 U10404 ( .A(n9958), .ZN(n9960) );
  NAND2_X2 U10405 ( .A1(n9960), .A2(n9959), .ZN(n9961) );
  NAND2_X2 U10406 ( .A1(n9962), .A2(n9961), .ZN(n9963) );
  AOI21_X4 U10407 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n9984) );
  INV_X4 U10408 ( .A(pipeline_alu_src_a[19]), .ZN(n11548) );
  OAI22_X2 U10409 ( .A1(n9447), .A2(n7134), .B1(n9966), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[19]) );
  INV_X4 U10410 ( .A(pipeline_rs2_data_bypassed[19]), .ZN(n9968) );
  OAI221_X2 U10411 ( .B1(n9968), .B2(n10056), .C1(n9270), .C2(n9396), .A(n9967), .ZN(pipeline_alu_src_b[19]) );
  INV_X4 U10412 ( .A(pipeline_alu_src_b[19]), .ZN(n9969) );
  OAI22_X2 U10413 ( .A1(n11548), .A2(n9453), .B1(n9969), .B2(n6744), .ZN(n9976) );
  OAI22_X2 U10414 ( .A1(n9969), .A2(n9453), .B1(n11548), .B2(n6744), .ZN(n9981) );
  INV_X4 U10415 ( .A(n9981), .ZN(n9970) );
  NAND2_X2 U10416 ( .A1(n9976), .A2(n9970), .ZN(n9975) );
  INV_X4 U10417 ( .A(n9971), .ZN(n9972) );
  NAND2_X2 U10418 ( .A1(n9973), .A2(n9972), .ZN(n9974) );
  NAND2_X2 U10419 ( .A1(n9975), .A2(n9974), .ZN(n9983) );
  INV_X4 U10420 ( .A(n9976), .ZN(n9980) );
  INV_X4 U10421 ( .A(n9977), .ZN(n9978) );
  OAI21_X4 U10422 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(n9995) );
  OAI22_X2 U10423 ( .A1(n7061), .A2(n7133), .B1(n9985), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[22]) );
  INV_X4 U10424 ( .A(pipeline_rs2_data_bypassed[22]), .ZN(n9986) );
  OAI221_X2 U10425 ( .B1(n9986), .B2(n10056), .C1(n702), .C2(n9397), .A(n10043), .ZN(pipeline_alu_src_b[22]) );
  INV_X4 U10426 ( .A(pipeline_alu_src_b[22]), .ZN(n9987) );
  OAI22_X2 U10427 ( .A1(n9987), .A2(n9456), .B1(n6624), .B2(n9451), .ZN(n10001) );
  OAI22_X2 U10428 ( .A1(n6624), .A2(n9453), .B1(n9987), .B2(n9451), .ZN(n10003) );
  INV_X4 U10429 ( .A(n10003), .ZN(n9988) );
  NAND2_X2 U10430 ( .A1(n10001), .A2(n9988), .ZN(n9993) );
  INV_X4 U10431 ( .A(n9989), .ZN(n9990) );
  NAND2_X2 U10432 ( .A1(n9991), .A2(n9990), .ZN(n9992) );
  NAND2_X2 U10433 ( .A1(n9993), .A2(n9992), .ZN(n9994) );
  INV_X4 U10434 ( .A(n6980), .ZN(n11847) );
  OAI22_X2 U10435 ( .A1(n7061), .A2(n7123), .B1(n9997), .B2(n10055), .ZN(
        pipeline_rs2_data_bypassed[23]) );
  INV_X4 U10436 ( .A(pipeline_rs2_data_bypassed[23]), .ZN(n9998) );
  OAI221_X2 U10437 ( .B1(n9998), .B2(n9448), .C1(n8223), .C2(n10044), .A(
        n10043), .ZN(pipeline_alu_src_b[23]) );
  INV_X4 U10438 ( .A(pipeline_alu_src_b[23]), .ZN(n9999) );
  OAI22_X2 U10439 ( .A1(n11847), .A2(n9453), .B1(n9999), .B2(n9451), .ZN(
        n10006) );
  OAI22_X2 U10440 ( .A1(n9999), .A2(n9453), .B1(n11847), .B2(n9451), .ZN(
        n10011) );
  INV_X4 U10441 ( .A(n10011), .ZN(n10000) );
  NAND2_X2 U10442 ( .A1(n10006), .A2(n10000), .ZN(n10005) );
  INV_X4 U10443 ( .A(n10001), .ZN(n10002) );
  NAND2_X2 U10444 ( .A1(n10003), .A2(n10002), .ZN(n10004) );
  NAND2_X2 U10445 ( .A1(n10005), .A2(n10004), .ZN(n10013) );
  INV_X4 U10446 ( .A(n10006), .ZN(n10010) );
  INV_X4 U10447 ( .A(n10007), .ZN(n10008) );
  INV_X4 U10448 ( .A(pipeline_rs2_data_bypassed[26]), .ZN(n10015) );
  OAI221_X2 U10449 ( .B1(n10015), .B2(n9448), .C1(n10338), .C2(n9396), .A(
        n10043), .ZN(pipeline_alu_src_b[26]) );
  INV_X4 U10450 ( .A(n6560), .ZN(n12099) );
  OAI22_X2 U10451 ( .A1(n10016), .A2(n9456), .B1(n12099), .B2(n9451), .ZN(
        n10029) );
  OAI22_X2 U10452 ( .A1(n12099), .A2(n9453), .B1(n10016), .B2(n9451), .ZN(
        n10031) );
  INV_X4 U10453 ( .A(n10031), .ZN(n10017) );
  NAND2_X2 U10454 ( .A1(n10029), .A2(n10017), .ZN(n10022) );
  INV_X4 U10455 ( .A(n10018), .ZN(n10019) );
  NAND2_X2 U10456 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  NAND2_X2 U10457 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  INV_X4 U10458 ( .A(pipeline_rs2_data_bypassed[27]), .ZN(n10026) );
  OAI22_X2 U10459 ( .A1(n6601), .A2(n9453), .B1(n10027), .B2(n9451), .ZN(
        n10034) );
  OAI22_X2 U10460 ( .A1(n10027), .A2(n9453), .B1(n6601), .B2(n9451), .ZN(
        n10039) );
  INV_X4 U10461 ( .A(n10039), .ZN(n10028) );
  NAND2_X2 U10462 ( .A1(n10034), .A2(n10028), .ZN(n10033) );
  INV_X4 U10463 ( .A(n10029), .ZN(n10030) );
  NAND2_X2 U10464 ( .A1(n10031), .A2(n10030), .ZN(n10032) );
  NAND2_X2 U10465 ( .A1(n10033), .A2(n10032), .ZN(n10041) );
  INV_X4 U10466 ( .A(n10034), .ZN(n10038) );
  INV_X4 U10467 ( .A(n10035), .ZN(n10036) );
  OAI22_X2 U10468 ( .A1(n12854), .A2(n10055), .B1(n9447), .B2(n7137), .ZN(
        pipeline_rs2_data_bypassed[30]) );
  INV_X4 U10469 ( .A(pipeline_rs2_data_bypassed[30]), .ZN(n10045) );
  INV_X4 U10470 ( .A(pipeline_alu_src_b[30]), .ZN(n12638) );
  OAI22_X2 U10471 ( .A1(n12638), .A2(n9456), .B1(n12635), .B2(n9451), .ZN(
        n10059) );
  OAI22_X2 U10472 ( .A1(n12635), .A2(n9453), .B1(n12638), .B2(n9451), .ZN(
        n10061) );
  INV_X4 U10473 ( .A(n10061), .ZN(n10046) );
  NAND2_X2 U10474 ( .A1(n10059), .A2(n10046), .ZN(n10051) );
  INV_X4 U10475 ( .A(n10047), .ZN(n10048) );
  NAND2_X2 U10476 ( .A1(n10049), .A2(n10048), .ZN(n10050) );
  NAND2_X2 U10477 ( .A1(n10051), .A2(n10050), .ZN(n10052) );
  INV_X4 U10478 ( .A(n7005), .ZN(n12593) );
  OAI22_X2 U10479 ( .A1(n12852), .A2(n10055), .B1(n9447), .B2(n7143), .ZN(
        pipeline_rs2_data_bypassed[31]) );
  INV_X4 U10480 ( .A(pipeline_rs2_data_bypassed[31]), .ZN(n12686) );
  OAI22_X2 U10481 ( .A1(n12593), .A2(n9453), .B1(n12566), .B2(n9451), .ZN(
        n10065) );
  INV_X4 U10482 ( .A(n10065), .ZN(n10058) );
  OAI22_X2 U10483 ( .A1(n12566), .A2(n9454), .B1(n12593), .B2(n9451), .ZN(
        n10064) );
  NAND2_X2 U10484 ( .A1(n10058), .A2(n10064), .ZN(n10063) );
  INV_X4 U10485 ( .A(n10059), .ZN(n10060) );
  NAND2_X2 U10486 ( .A1(n10061), .A2(n10060), .ZN(n10062) );
  NAND2_X2 U10487 ( .A1(n10063), .A2(n10062), .ZN(n10068) );
  INV_X4 U10488 ( .A(n10064), .ZN(n10066) );
  NAND2_X2 U10489 ( .A1(n10066), .A2(n10065), .ZN(n10067) );
  NAND3_X2 U10490 ( .A1(n10081), .A2(n6578), .A3(n10085), .ZN(n12357) );
  NOR2_X2 U10491 ( .A1(n6617), .A2(n12357), .ZN(n10070) );
  NAND2_X2 U10492 ( .A1(n12793), .A2(n10081), .ZN(n12783) );
  NOR2_X2 U10493 ( .A1(n10070), .A2(n9513), .ZN(n10071) );
  NOR2_X2 U10494 ( .A1(n6943), .A2(n10071), .ZN(n10079) );
  MUX2_X2 U10495 ( .A(pipeline_alu_N320), .B(pipeline_alu_N319), .S(n10081), 
        .Z(n10072) );
  NAND2_X2 U10496 ( .A1(n10072), .A2(n10083), .ZN(n10076) );
  MUX2_X2 U10497 ( .A(pipeline_alu_N252), .B(pipeline_alu_N251), .S(n10081), 
        .Z(n10073) );
  NAND2_X2 U10498 ( .A1(n10074), .A2(n10073), .ZN(n10075) );
  MUX2_X2 U10499 ( .A(n12793), .B(n9479), .S(n6943), .Z(n10084) );
  NOR2_X2 U10500 ( .A1(n9513), .A2(n10084), .ZN(n10086) );
  NAND2_X2 U10501 ( .A1(n7068), .A2(n10085), .ZN(n12590) );
  INV_X4 U10502 ( .A(n12590), .ZN(n12662) );
  OAI22_X2 U10503 ( .A1(n11404), .A2(n10086), .B1(n12785), .B2(n11372), .ZN(
        n10087) );
  AOI221_X2 U10504 ( .B1(pipeline_alu_N253), .B2(n6812), .C1(pipeline_alu_N59), 
        .C2(n6813), .A(n10087), .ZN(n10088) );
  NAND2_X2 U10505 ( .A1(n10089), .A2(n10088), .ZN(dmem_haddr[0]) );
  NAND3_X2 U10506 ( .A1(n13097), .A2(n12402), .A3(dmem_haddr[0]), .ZN(n10090)
         );
  NAND2_X2 U10507 ( .A1(n10091), .A2(n10090), .ZN(n10304) );
  INV_X4 U10508 ( .A(n10304), .ZN(n11178) );
  NAND2_X2 U10509 ( .A1(n11178), .A2(n6799), .ZN(n10094) );
  NOR3_X2 U10510 ( .A1(n10094), .A2(n10093), .A3(n10385), .ZN(n10095) );
  NAND3_X2 U10511 ( .A1(n6922), .A2(n10096), .A3(n10095), .ZN(n10388) );
  NAND2_X2 U10512 ( .A1(n12832), .A2(n10388), .ZN(n10345) );
  NAND2_X2 U10513 ( .A1(n10345), .A2(n13130), .ZN(n12831) );
  AOI221_X2 U10514 ( .B1(imem_hrdata[4]), .B2(n12832), .C1(n9517), .C2(
        pipeline_inst_DX[4]), .A(n12831), .ZN(n10097) );
  INV_X4 U10515 ( .A(n10097), .ZN(n6259) );
  INV_X4 U10516 ( .A(imem_hrdata[2]), .ZN(n10099) );
  OAI22_X2 U10517 ( .A1(n6639), .A2(n10099), .B1(n9623), .B2(n12823), .ZN(
        n6257) );
  INV_X4 U10518 ( .A(imem_hrdata[5]), .ZN(n10100) );
  OAI22_X2 U10519 ( .A1(n6639), .A2(n10100), .B1(n9651), .B2(n12823), .ZN(
        n6260) );
  INV_X4 U10520 ( .A(imem_hrdata[6]), .ZN(n10101) );
  OAI22_X2 U10521 ( .A1(n6639), .A2(n10101), .B1(n9650), .B2(n12823), .ZN(
        n6261) );
  INV_X4 U10522 ( .A(imem_hrdata[3]), .ZN(n10102) );
  OAI22_X2 U10523 ( .A1(n6639), .A2(n10102), .B1(n9648), .B2(n12823), .ZN(
        n6258) );
  INV_X4 U10524 ( .A(imem_hrdata[31]), .ZN(n10103) );
  OAI22_X2 U10525 ( .A1(n6639), .A2(n10103), .B1(n10242), .B2(n12823), .ZN(
        n6295) );
  INV_X4 U10526 ( .A(imem_hrdata[30]), .ZN(n10104) );
  INV_X4 U10527 ( .A(imem_hrdata[7]), .ZN(n10105) );
  INV_X4 U10528 ( .A(imem_hrdata[8]), .ZN(n10106) );
  INV_X4 U10529 ( .A(imem_hrdata[9]), .ZN(n10107) );
  INV_X4 U10530 ( .A(imem_hrdata[17]), .ZN(n10108) );
  INV_X4 U10531 ( .A(imem_hrdata[18]), .ZN(n10109) );
  INV_X4 U10532 ( .A(imem_hrdata[19]), .ZN(n10110) );
  INV_X4 U10533 ( .A(imem_hrdata[16]), .ZN(n10111) );
  INV_X4 U10534 ( .A(imem_hrdata[15]), .ZN(n10112) );
  INV_X4 U10535 ( .A(imem_hrdata[11]), .ZN(n10113) );
  INV_X4 U10536 ( .A(imem_hrdata[10]), .ZN(n10114) );
  INV_X4 U10537 ( .A(imem_hrdata[14]), .ZN(n10115) );
  INV_X4 U10538 ( .A(imem_hrdata[12]), .ZN(n10116) );
  OAI22_X2 U10539 ( .A1(n6639), .A2(n10116), .B1(n601), .B2(n12823), .ZN(n6273) );
  INV_X4 U10540 ( .A(imem_hrdata[13]), .ZN(n10117) );
  INV_X4 U10541 ( .A(imem_hrdata[22]), .ZN(n10118) );
  OAI22_X2 U10542 ( .A1(n6639), .A2(n10118), .B1(n702), .B2(n12823), .ZN(n6285) );
  INV_X4 U10543 ( .A(imem_hrdata[24]), .ZN(n10119) );
  OAI22_X2 U10544 ( .A1(n6639), .A2(n10119), .B1(n8214), .B2(n12823), .ZN(
        n6287) );
  INV_X4 U10545 ( .A(imem_hrdata[25]), .ZN(n10120) );
  OAI22_X2 U10546 ( .A1(n6639), .A2(n10120), .B1(n10336), .B2(n12823), .ZN(
        n6288) );
  INV_X4 U10547 ( .A(imem_hrdata[27]), .ZN(n10121) );
  INV_X4 U10548 ( .A(imem_hrdata[26]), .ZN(n10122) );
  INV_X4 U10549 ( .A(imem_hrdata[29]), .ZN(n10123) );
  OAI22_X2 U10550 ( .A1(n6639), .A2(n10123), .B1(n9632), .B2(n12823), .ZN(
        n6292) );
  INV_X4 U10551 ( .A(imem_hrdata[23]), .ZN(n10124) );
  OAI22_X2 U10552 ( .A1(n6639), .A2(n10124), .B1(n8223), .B2(n12823), .ZN(
        n6286) );
  INV_X4 U10553 ( .A(imem_hrdata[28]), .ZN(n10125) );
  OAI22_X2 U10554 ( .A1(n6639), .A2(n10125), .B1(n9634), .B2(n12823), .ZN(
        n6291) );
  INV_X4 U10555 ( .A(imem_hrdata[20]), .ZN(n10126) );
  NOR2_X2 U10556 ( .A1(n10127), .A2(n12827), .ZN(n6299) );
  NAND3_X2 U10557 ( .A1(n10130), .A2(n10129), .A3(n10128), .ZN(n10135) );
  NOR2_X2 U10558 ( .A1(n10132), .A2(n10131), .ZN(n10133) );
  NOR3_X2 U10559 ( .A1(n10135), .A2(n10134), .A3(n10133), .ZN(n10136) );
  NAND2_X2 U10560 ( .A1(n9525), .A2(n13097), .ZN(n12826) );
  NAND2_X2 U10561 ( .A1(n12827), .A2(n13130), .ZN(n12829) );
  OAI22_X2 U10562 ( .A1(n10136), .A2(n12826), .B1(n791), .B2(n12829), .ZN(
        n6252) );
  MUX2_X2 U10563 ( .A(n12992), .B(pipeline_inst_DX[11]), .S(n9525), .Z(n6270)
         );
  MUX2_X2 U10564 ( .A(n12995), .B(pipeline_inst_DX[10]), .S(n9524), .Z(n6268)
         );
  MUX2_X2 U10565 ( .A(pipeline_reg_to_wr_WB[1]), .B(n10137), .S(n9522), .Z(
        n6264) );
  MUX2_X2 U10566 ( .A(pipeline_reg_to_wr_WB[2]), .B(pipeline_inst_DX[9]), .S(
        n9523), .Z(n6266) );
  MUX2_X2 U10567 ( .A(n12990), .B(n10138), .S(n9525), .Z(n6262) );
  NAND2_X2 U10568 ( .A1(n10139), .A2(n13097), .ZN(n13125) );
  OAI22_X2 U10569 ( .A1(n790), .A2(n12829), .B1(n12827), .B2(n13125), .ZN(
        n6253) );
  NAND2_X2 U10570 ( .A1(n12835), .A2(n13097), .ZN(n10140) );
  NAND2_X2 U10571 ( .A1(n10140), .A2(n13125), .ZN(dmem_htrans[1]) );
  INV_X4 U10572 ( .A(dmem_htrans[1]), .ZN(n10141) );
  OAI22_X2 U10573 ( .A1(n789), .A2(n12829), .B1(n10141), .B2(n12827), .ZN(
        n6254) );
  NAND2_X2 U10574 ( .A1(n12834), .A2(n13096), .ZN(n10142) );
  NAND2_X2 U10575 ( .A1(n10142), .A2(n12836), .ZN(n10143) );
  MUX2_X2 U10576 ( .A(n10144), .B(n10143), .S(n9525), .Z(n6333) );
  NAND2_X2 U10577 ( .A1(n9642), .A2(pipeline_md_state[0]), .ZN(n13029) );
  NOR2_X2 U10578 ( .A1(n1558), .A2(n9518), .ZN(n10145) );
  NAND2_X2 U10579 ( .A1(n13097), .A2(n7085), .ZN(n12828) );
  INV_X4 U10580 ( .A(n12828), .ZN(n10195) );
  NAND2_X2 U10581 ( .A1(n6810), .A2(pipeline_md_state[1]), .ZN(n10200) );
  INV_X4 U10582 ( .A(n10200), .ZN(n10269) );
  NOR3_X2 U10583 ( .A1(n10145), .A2(n10195), .A3(n10269), .ZN(n10146) );
  NOR2_X2 U10584 ( .A1(htif_reset), .A2(n10146), .ZN(pipeline_md_N161) );
  INV_X4 U10585 ( .A(n1558), .ZN(n10147) );
  NOR2_X2 U10586 ( .A1(n9518), .A2(n10147), .ZN(n10148) );
  NOR2_X2 U10587 ( .A1(n10269), .A2(n10148), .ZN(n10149) );
  NOR2_X2 U10588 ( .A1(htif_reset), .A2(n10149), .ZN(pipeline_md_N162) );
  MUX2_X2 U10589 ( .A(n10150), .B(n10193), .S(n10195), .Z(n6242) );
  NOR2_X2 U10590 ( .A1(dmem_hsize[1]), .A2(n603), .ZN(n10151) );
  MUX2_X2 U10591 ( .A(pipeline_md_op_0_), .B(n10151), .S(n10195), .Z(n6243) );
  NAND2_X2 U10592 ( .A1(n964), .A2(n963), .ZN(n10197) );
  NAND2_X2 U10593 ( .A1(n9519), .A2(n10197), .ZN(n10201) );
  INV_X4 U10594 ( .A(n10201), .ZN(n10271) );
  NAND2_X2 U10595 ( .A1(pipeline_md_a_geq), .A2(n10271), .ZN(n10152) );
  NAND2_X2 U10596 ( .A1(n10152), .A2(n12828), .ZN(n12763) );
  NAND2_X2 U10597 ( .A1(n9519), .A2(n9504), .ZN(n12765) );
  INV_X4 U10598 ( .A(pipeline_md_N313), .ZN(n10153) );
  OAI22_X2 U10599 ( .A1(n9505), .A2(n10153), .B1(n1149), .B2(n12763), .ZN(
        n5715) );
  INV_X4 U10600 ( .A(pipeline_md_N312), .ZN(n10154) );
  OAI22_X2 U10601 ( .A1(n9505), .A2(n10154), .B1(n1148), .B2(n12763), .ZN(
        n5714) );
  INV_X4 U10602 ( .A(pipeline_md_N311), .ZN(n10155) );
  OAI22_X2 U10603 ( .A1(n9505), .A2(n10155), .B1(n1147), .B2(n12763), .ZN(
        n5713) );
  INV_X4 U10604 ( .A(pipeline_md_N310), .ZN(n10156) );
  OAI22_X2 U10605 ( .A1(n9505), .A2(n10156), .B1(n1146), .B2(n12763), .ZN(
        n5712) );
  INV_X4 U10606 ( .A(pipeline_md_N309), .ZN(n10157) );
  OAI22_X2 U10607 ( .A1(n9505), .A2(n10157), .B1(n1145), .B2(n12763), .ZN(
        n5711) );
  INV_X4 U10608 ( .A(pipeline_md_N308), .ZN(n10158) );
  OAI22_X2 U10609 ( .A1(n9505), .A2(n10158), .B1(n1144), .B2(n12763), .ZN(
        n5710) );
  INV_X4 U10610 ( .A(pipeline_md_N307), .ZN(n10159) );
  INV_X4 U10612 ( .A(pipeline_md_N306), .ZN(n10160) );
  INV_X4 U10614 ( .A(pipeline_md_N305), .ZN(n10161) );
  INV_X4 U10616 ( .A(pipeline_md_N304), .ZN(n10162) );
  INV_X4 U10618 ( .A(pipeline_md_N303), .ZN(n10163) );
  OAI22_X2 U10619 ( .A1(n9505), .A2(n10163), .B1(n1139), .B2(n9504), .ZN(n5705) );
  INV_X4 U10620 ( .A(pipeline_md_N302), .ZN(n10164) );
  OAI22_X2 U10621 ( .A1(n9505), .A2(n10164), .B1(n1138), .B2(n9504), .ZN(n5704) );
  INV_X4 U10622 ( .A(pipeline_md_N301), .ZN(n10165) );
  OAI22_X2 U10623 ( .A1(n9505), .A2(n10165), .B1(n1137), .B2(n9504), .ZN(n5703) );
  INV_X4 U10624 ( .A(pipeline_md_N300), .ZN(n10166) );
  OAI22_X2 U10625 ( .A1(n9505), .A2(n10166), .B1(n1136), .B2(n9504), .ZN(n5702) );
  INV_X4 U10626 ( .A(pipeline_md_N299), .ZN(n10167) );
  OAI22_X2 U10627 ( .A1(n9505), .A2(n10167), .B1(n1135), .B2(n9504), .ZN(n5701) );
  INV_X4 U10628 ( .A(pipeline_md_N298), .ZN(n10168) );
  OAI22_X2 U10629 ( .A1(n9505), .A2(n10168), .B1(n1134), .B2(n9504), .ZN(n5700) );
  INV_X4 U10630 ( .A(pipeline_md_N297), .ZN(n10169) );
  OAI22_X2 U10631 ( .A1(n9505), .A2(n10169), .B1(n1133), .B2(n9504), .ZN(n5699) );
  INV_X4 U10632 ( .A(pipeline_md_N296), .ZN(n10170) );
  OAI22_X2 U10633 ( .A1(n9505), .A2(n10170), .B1(n1132), .B2(n9504), .ZN(n5698) );
  INV_X4 U10634 ( .A(pipeline_md_N295), .ZN(n10171) );
  OAI22_X2 U10635 ( .A1(n9505), .A2(n10171), .B1(n1131), .B2(n9504), .ZN(n5697) );
  INV_X4 U10636 ( .A(pipeline_md_N294), .ZN(n10172) );
  OAI22_X2 U10637 ( .A1(n9505), .A2(n10172), .B1(n1130), .B2(n9504), .ZN(n5696) );
  INV_X4 U10638 ( .A(pipeline_md_N293), .ZN(n10173) );
  OAI22_X2 U10639 ( .A1(n9505), .A2(n10173), .B1(n1129), .B2(n9504), .ZN(n5695) );
  INV_X4 U10640 ( .A(pipeline_md_N292), .ZN(n10174) );
  OAI22_X2 U10641 ( .A1(n9505), .A2(n10174), .B1(n1128), .B2(n9504), .ZN(n5694) );
  INV_X4 U10642 ( .A(pipeline_md_N291), .ZN(n10175) );
  OAI22_X2 U10643 ( .A1(n9505), .A2(n10175), .B1(n1127), .B2(n9504), .ZN(n5693) );
  INV_X4 U10644 ( .A(pipeline_md_N290), .ZN(n10176) );
  OAI22_X2 U10645 ( .A1(n9505), .A2(n10176), .B1(n1126), .B2(n9504), .ZN(n5692) );
  INV_X4 U10646 ( .A(pipeline_md_N289), .ZN(n10177) );
  OAI22_X2 U10647 ( .A1(n9505), .A2(n10177), .B1(n1125), .B2(n9504), .ZN(n5691) );
  INV_X4 U10648 ( .A(pipeline_md_N288), .ZN(n10178) );
  OAI22_X2 U10649 ( .A1(n9505), .A2(n10178), .B1(n1124), .B2(n9504), .ZN(n5690) );
  INV_X4 U10650 ( .A(pipeline_md_N287), .ZN(n10179) );
  OAI22_X2 U10651 ( .A1(n9505), .A2(n10179), .B1(n1123), .B2(n9504), .ZN(n5689) );
  INV_X4 U10652 ( .A(pipeline_md_N286), .ZN(n10180) );
  OAI22_X2 U10653 ( .A1(n9505), .A2(n10180), .B1(n1122), .B2(n12763), .ZN(
        n5688) );
  INV_X4 U10654 ( .A(pipeline_md_N285), .ZN(n10181) );
  OAI22_X2 U10655 ( .A1(n9505), .A2(n10181), .B1(n1121), .B2(n12763), .ZN(
        n5687) );
  INV_X4 U10656 ( .A(pipeline_md_N284), .ZN(n10182) );
  OAI22_X2 U10657 ( .A1(n9505), .A2(n10182), .B1(n1120), .B2(n12763), .ZN(
        n5686) );
  INV_X4 U10658 ( .A(pipeline_md_N283), .ZN(n10183) );
  OAI22_X2 U10659 ( .A1(n9505), .A2(n10183), .B1(n1119), .B2(n12763), .ZN(
        n5685) );
  NAND3_X2 U10660 ( .A1(n10186), .A2(n10185), .A3(n10184), .ZN(n10188) );
  NAND2_X2 U10661 ( .A1(n10187), .A2(pipeline_rs1_data_bypassed[31]), .ZN(
        n10265) );
  INV_X4 U10662 ( .A(n10265), .ZN(n10264) );
  NOR2_X2 U10663 ( .A1(pipeline_md_op_0_), .A2(n964), .ZN(n10189) );
  NAND2_X2 U10664 ( .A1(n10188), .A2(pipeline_rs2_data_bypassed[31]), .ZN(
        n12683) );
  NOR2_X2 U10665 ( .A1(n10189), .A2(n12683), .ZN(n10190) );
  XOR2_X2 U10666 ( .A(n10264), .B(n10190), .Z(n10191) );
  MUX2_X2 U10667 ( .A(n10192), .B(n10191), .S(n10195), .Z(n6241) );
  MUX2_X2 U10668 ( .A(pipeline_md_out_sel[1]), .B(n10193), .S(n10195), .Z(
        n6244) );
  NOR2_X2 U10669 ( .A1(n10194), .A2(pipeline_dmem_type_2_), .ZN(n10196) );
  MUX2_X2 U10670 ( .A(pipeline_md_out_sel[0]), .B(n10196), .S(n10195), .Z(
        n6245) );
  INV_X4 U10671 ( .A(n10197), .ZN(n10198) );
  NAND2_X2 U10672 ( .A1(pipeline_md_N185), .A2(n6918), .ZN(n10199) );
  NAND3_X2 U10673 ( .A1(n9503), .A2(n10200), .A3(n10199), .ZN(n10277) );
  NAND2_X2 U10674 ( .A1(n6918), .A2(n10277), .ZN(n12753) );
  INV_X4 U10675 ( .A(pipeline_md_N248), .ZN(n10202) );
  OAI22_X2 U10676 ( .A1(n9501), .A2(n10202), .B1(n958), .B2(n6809), .ZN(n5591)
         );
  INV_X4 U10677 ( .A(pipeline_md_N247), .ZN(n10203) );
  OAI22_X2 U10678 ( .A1(n9501), .A2(n10203), .B1(n956), .B2(n6809), .ZN(n5592)
         );
  INV_X4 U10679 ( .A(pipeline_md_N246), .ZN(n10204) );
  OAI22_X2 U10680 ( .A1(n9501), .A2(n10204), .B1(n954), .B2(n6809), .ZN(n5593)
         );
  INV_X4 U10681 ( .A(pipeline_md_N245), .ZN(n10205) );
  OAI22_X2 U10682 ( .A1(n9501), .A2(n10205), .B1(n952), .B2(n6809), .ZN(n5594)
         );
  INV_X4 U10683 ( .A(pipeline_md_N244), .ZN(n10206) );
  OAI22_X2 U10684 ( .A1(n9501), .A2(n10206), .B1(n950), .B2(n6809), .ZN(n5595)
         );
  INV_X4 U10685 ( .A(pipeline_md_N243), .ZN(n10207) );
  INV_X4 U10687 ( .A(pipeline_md_N242), .ZN(n10208) );
  INV_X4 U10689 ( .A(pipeline_md_N241), .ZN(n10209) );
  INV_X4 U10691 ( .A(pipeline_md_N240), .ZN(n10210) );
  INV_X4 U10693 ( .A(pipeline_md_N239), .ZN(n10211) );
  INV_X4 U10695 ( .A(pipeline_md_N238), .ZN(n10212) );
  INV_X4 U10697 ( .A(pipeline_md_N237), .ZN(n10213) );
  INV_X4 U10699 ( .A(pipeline_md_N236), .ZN(n10214) );
  OAI22_X2 U10700 ( .A1(n12753), .A2(n10214), .B1(n934), .B2(n6809), .ZN(n5603) );
  INV_X4 U10701 ( .A(pipeline_md_N235), .ZN(n10215) );
  OAI22_X2 U10702 ( .A1(n12753), .A2(n10215), .B1(n932), .B2(n6809), .ZN(n5604) );
  INV_X4 U10703 ( .A(pipeline_md_N234), .ZN(n10216) );
  OAI22_X2 U10704 ( .A1(n12753), .A2(n10216), .B1(n930), .B2(n6809), .ZN(n5605) );
  INV_X4 U10705 ( .A(pipeline_md_N233), .ZN(n10217) );
  OAI22_X2 U10706 ( .A1(n12753), .A2(n10217), .B1(n928), .B2(n6809), .ZN(n5606) );
  INV_X4 U10707 ( .A(pipeline_md_N232), .ZN(n10218) );
  OAI22_X2 U10708 ( .A1(n12753), .A2(n10218), .B1(n926), .B2(n6809), .ZN(n5607) );
  INV_X4 U10709 ( .A(pipeline_md_N231), .ZN(n10219) );
  OAI22_X2 U10710 ( .A1(n12753), .A2(n10219), .B1(n924), .B2(n6809), .ZN(n5608) );
  INV_X4 U10711 ( .A(pipeline_md_N230), .ZN(n10220) );
  OAI22_X2 U10712 ( .A1(n12753), .A2(n10220), .B1(n922), .B2(n6809), .ZN(n5609) );
  INV_X4 U10713 ( .A(pipeline_md_N229), .ZN(n10221) );
  OAI22_X2 U10714 ( .A1(n12753), .A2(n10221), .B1(n920), .B2(n6809), .ZN(n5610) );
  INV_X4 U10715 ( .A(pipeline_md_N228), .ZN(n10222) );
  OAI22_X2 U10716 ( .A1(n12753), .A2(n10222), .B1(n918), .B2(n6809), .ZN(n5611) );
  INV_X4 U10717 ( .A(pipeline_md_N227), .ZN(n10223) );
  OAI22_X2 U10718 ( .A1(n12753), .A2(n10223), .B1(n916), .B2(n6809), .ZN(n5612) );
  INV_X4 U10719 ( .A(pipeline_md_N226), .ZN(n10224) );
  OAI22_X2 U10720 ( .A1(n12753), .A2(n10224), .B1(n914), .B2(n6809), .ZN(n5613) );
  INV_X4 U10721 ( .A(pipeline_md_N225), .ZN(n10225) );
  OAI22_X2 U10722 ( .A1(n12753), .A2(n10225), .B1(n912), .B2(n6809), .ZN(n5614) );
  INV_X4 U10723 ( .A(pipeline_md_N224), .ZN(n10226) );
  OAI22_X2 U10724 ( .A1(n12753), .A2(n10226), .B1(n910), .B2(n6809), .ZN(n5615) );
  INV_X4 U10725 ( .A(pipeline_md_N223), .ZN(n10227) );
  OAI22_X2 U10726 ( .A1(n12753), .A2(n10227), .B1(n908), .B2(n6809), .ZN(n5616) );
  INV_X4 U10727 ( .A(pipeline_md_N222), .ZN(n10228) );
  OAI22_X2 U10728 ( .A1(n12753), .A2(n10228), .B1(n906), .B2(n6809), .ZN(n5617) );
  INV_X4 U10729 ( .A(pipeline_md_N221), .ZN(n10229) );
  OAI22_X2 U10730 ( .A1(n12753), .A2(n10229), .B1(n904), .B2(n6809), .ZN(n5618) );
  INV_X4 U10731 ( .A(pipeline_md_N220), .ZN(n10230) );
  OAI22_X2 U10732 ( .A1(n12753), .A2(n10230), .B1(n902), .B2(n6809), .ZN(n5619) );
  INV_X4 U10733 ( .A(pipeline_md_N219), .ZN(n10231) );
  OAI22_X2 U10734 ( .A1(n12753), .A2(n10231), .B1(n900), .B2(n6809), .ZN(n5620) );
  INV_X4 U10735 ( .A(pipeline_md_N218), .ZN(n10232) );
  OAI22_X2 U10736 ( .A1(n9501), .A2(n10232), .B1(n898), .B2(n6809), .ZN(n5621)
         );
  NAND2_X2 U10737 ( .A1(pipeline_md_out_sel[1]), .A2(n1153), .ZN(n10276) );
  MUX2_X2 U10738 ( .A(n10234), .B(n10233), .S(n9499), .Z(
        pipeline_md_result_muxed[63]) );
  MUX2_X2 U10739 ( .A(pipeline_md_result[62]), .B(pipeline_md_a[62]), .S(n9500), .Z(pipeline_md_result_muxed[62]) );
  MUX2_X2 U10740 ( .A(pipeline_md_result[61]), .B(pipeline_md_a[61]), .S(n9499), .Z(pipeline_md_result_muxed[61]) );
  MUX2_X2 U10741 ( .A(pipeline_md_result[60]), .B(pipeline_md_a[60]), .S(n9500), .Z(pipeline_md_result_muxed[60]) );
  MUX2_X2 U10742 ( .A(pipeline_md_result[59]), .B(pipeline_md_a[59]), .S(n9499), .Z(pipeline_md_result_muxed[59]) );
  MUX2_X2 U10743 ( .A(pipeline_md_result[58]), .B(pipeline_md_a[58]), .S(n9500), .Z(pipeline_md_result_muxed[58]) );
  MUX2_X2 U10744 ( .A(pipeline_md_result[57]), .B(pipeline_md_a[57]), .S(n9499), .Z(pipeline_md_result_muxed[57]) );
  MUX2_X2 U10745 ( .A(pipeline_md_result[56]), .B(pipeline_md_a[56]), .S(n9500), .Z(pipeline_md_result_muxed[56]) );
  MUX2_X2 U10746 ( .A(pipeline_md_result[55]), .B(pipeline_md_a[55]), .S(n9499), .Z(pipeline_md_result_muxed[55]) );
  MUX2_X2 U10747 ( .A(pipeline_md_result[54]), .B(pipeline_md_a[54]), .S(n9500), .Z(pipeline_md_result_muxed[54]) );
  MUX2_X2 U10748 ( .A(pipeline_md_result[53]), .B(pipeline_md_a[53]), .S(n9499), .Z(pipeline_md_result_muxed[53]) );
  MUX2_X2 U10749 ( .A(pipeline_md_result[52]), .B(pipeline_md_a[52]), .S(n9500), .Z(pipeline_md_result_muxed[52]) );
  MUX2_X2 U10750 ( .A(pipeline_md_result[51]), .B(pipeline_md_a[51]), .S(n9499), .Z(pipeline_md_result_muxed[51]) );
  MUX2_X2 U10751 ( .A(pipeline_md_result[50]), .B(pipeline_md_a[50]), .S(n9500), .Z(pipeline_md_result_muxed[50]) );
  MUX2_X2 U10752 ( .A(pipeline_md_result[49]), .B(pipeline_md_a[49]), .S(n9499), .Z(pipeline_md_result_muxed[49]) );
  MUX2_X2 U10753 ( .A(pipeline_md_result[48]), .B(pipeline_md_a[48]), .S(n9500), .Z(pipeline_md_result_muxed[48]) );
  MUX2_X2 U10754 ( .A(pipeline_md_result[47]), .B(pipeline_md_a[47]), .S(n9499), .Z(pipeline_md_result_muxed[47]) );
  MUX2_X2 U10755 ( .A(pipeline_md_result[46]), .B(pipeline_md_a[46]), .S(n9500), .Z(pipeline_md_result_muxed[46]) );
  MUX2_X2 U10756 ( .A(pipeline_md_result[45]), .B(pipeline_md_a[45]), .S(n9499), .Z(pipeline_md_result_muxed[45]) );
  MUX2_X2 U10757 ( .A(pipeline_md_result[44]), .B(pipeline_md_a[44]), .S(n9500), .Z(pipeline_md_result_muxed[44]) );
  MUX2_X2 U10758 ( .A(pipeline_md_result[43]), .B(pipeline_md_a[43]), .S(n9499), .Z(pipeline_md_result_muxed[43]) );
  MUX2_X2 U10759 ( .A(pipeline_md_result[42]), .B(pipeline_md_a[42]), .S(n9500), .Z(pipeline_md_result_muxed[42]) );
  MUX2_X2 U10760 ( .A(pipeline_md_result[41]), .B(pipeline_md_a[41]), .S(n9499), .Z(pipeline_md_result_muxed[41]) );
  MUX2_X2 U10761 ( .A(pipeline_md_result[40]), .B(pipeline_md_a[40]), .S(n9499), .Z(pipeline_md_result_muxed[40]) );
  MUX2_X2 U10762 ( .A(pipeline_md_result[39]), .B(pipeline_md_a[39]), .S(n9499), .Z(pipeline_md_result_muxed[39]) );
  MUX2_X2 U10763 ( .A(pipeline_md_result[38]), .B(pipeline_md_a[38]), .S(n9499), .Z(pipeline_md_result_muxed[38]) );
  MUX2_X2 U10764 ( .A(pipeline_md_result[37]), .B(pipeline_md_a[37]), .S(n9499), .Z(pipeline_md_result_muxed[37]) );
  MUX2_X2 U10765 ( .A(pipeline_md_result[36]), .B(pipeline_md_a[36]), .S(n9500), .Z(pipeline_md_result_muxed[36]) );
  MUX2_X2 U10766 ( .A(pipeline_md_result[35]), .B(pipeline_md_a[35]), .S(n9499), .Z(pipeline_md_result_muxed[35]) );
  MUX2_X2 U10767 ( .A(pipeline_md_result[34]), .B(pipeline_md_a[34]), .S(n9499), .Z(pipeline_md_result_muxed[34]) );
  MUX2_X2 U10768 ( .A(pipeline_md_result[33]), .B(pipeline_md_a[33]), .S(n9499), .Z(pipeline_md_result_muxed[33]) );
  MUX2_X2 U10769 ( .A(pipeline_md_result[32]), .B(pipeline_md_a[32]), .S(n9500), .Z(pipeline_md_result_muxed[32]) );
  MUX2_X2 U10770 ( .A(pipeline_md_resp_result[31]), .B(pipeline_md_a[31]), .S(
        n9500), .Z(pipeline_md_result_muxed[31]) );
  NAND2_X2 U10771 ( .A1(n7166), .A2(n7169), .ZN(n13103) );
  INV_X4 U10772 ( .A(n10237), .ZN(n10251) );
  NAND2_X2 U10773 ( .A1(n6641), .A2(n7077), .ZN(n13104) );
  NAND2_X2 U10774 ( .A1(n11229), .A2(n10238), .ZN(n10239) );
  OAI221_X2 U10775 ( .B1(n1545), .B2(n9462), .C1(n12665), .C2(n11262), .A(
        n10239), .ZN(n10240) );
  AOI221_X2 U10776 ( .B1(n11138), .B2(n10241), .C1(n11136), .C2(
        ext_interrupts[22]), .A(n10240), .ZN(n10257) );
  NAND3_X2 U10777 ( .A1(n7079), .A2(n7163), .A3(n10248), .ZN(n11261) );
  NAND2_X2 U10778 ( .A1(n7176), .A2(n7016), .ZN(n13111) );
  NAND3_X2 U10779 ( .A1(n6641), .A2(n6664), .A3(n7176), .ZN(n11269) );
  AOI221_X2 U10780 ( .B1(n9527), .B2(n10245), .C1(pipeline_csr_mtime_full[30]), 
        .C2(n13108), .A(n10244), .ZN(n10256) );
  NAND2_X2 U10781 ( .A1(n7166), .A2(n10248), .ZN(n13113) );
  NAND2_X2 U10782 ( .A1(pipeline_imm_31_), .A2(pipeline_inst_DX[30]), .ZN(
        n10247) );
  OAI33_X1 U10783 ( .A1(n10247), .A2(pipeline_inst_DX[28]), .A3(
        pipeline_inst_DX[29]), .B1(n10246), .B2(n9634), .B3(n10242), .ZN(
        n10339) );
  NAND2_X2 U10784 ( .A1(n7063), .A2(n9402), .ZN(n10783) );
  NAND3_X2 U10785 ( .A1(n7163), .A2(n7165), .A3(n7079), .ZN(n11235) );
  AOI221_X2 U10787 ( .B1(pipeline_csr_mscratch[30]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[30]), .C2(n13116), .A(n10250), .ZN(n10255) );
  OAI22_X2 U10788 ( .A1(n9460), .A2(n10252), .B1(n9526), .B2(n6830), .ZN(
        n10253) );
  AOI221_X2 U10789 ( .B1(pipeline_csr_instret_full[62]), .B2(n11105), .C1(
        pipeline_csr_time_full[62]), .C2(n11257), .A(n10253), .ZN(n10254) );
  NOR2_X2 U10790 ( .A1(pipeline_rs1_data_bypassed[30]), .A2(n9463), .ZN(n10259) );
  NOR2_X2 U10791 ( .A1(n6793), .A2(n10259), .ZN(n10262) );
  NAND2_X2 U10792 ( .A1(n7179), .A2(n7168), .ZN(n10260) );
  NAND2_X2 U10793 ( .A1(htif_pcr_req_data[30]), .A2(n13131), .ZN(n10261) );
  OAI221_X2 U10794 ( .B1(n7211), .B2(n10262), .C1(n12418), .C2(n9467), .A(
        n10261), .ZN(n12667) );
  INV_X4 U10795 ( .A(n12667), .ZN(n12670) );
  INV_X4 U10796 ( .A(n10341), .ZN(n10824) );
  NAND2_X2 U10797 ( .A1(n7192), .A2(n6843), .ZN(n10263) );
  OAI22_X2 U10798 ( .A1(n12670), .A2(n6690), .B1(n1221), .B2(n6708), .ZN(n6178) );
  OAI22_X2 U10799 ( .A1(n12670), .A2(n9516), .B1(n1545), .B2(n6660), .ZN(n6237) );
  INV_X4 U10800 ( .A(pipeline_md_N251), .ZN(n10266) );
  OAI22_X2 U10801 ( .A1(n1087), .A2(n9504), .B1(n9505), .B2(n10266), .ZN(
        n10267) );
  INV_X4 U10802 ( .A(n10268), .ZN(n5716) );
  NAND2_X2 U10803 ( .A1(pipeline_md_out_sel[0]), .A2(n1154), .ZN(n10275) );
  INV_X4 U10804 ( .A(n10275), .ZN(n10270) );
  INV_X4 U10805 ( .A(pipeline_md_result_muxed[32]), .ZN(n10273) );
  NOR2_X2 U10806 ( .A1(pipeline_md_N315), .A2(pipeline_md_resp_result[0]), 
        .ZN(n10272) );
  OAI22_X2 U10807 ( .A1(n10273), .A2(n6692), .B1(n10272), .B2(n6667), .ZN(
        n10274) );
  AOI221_X2 U10808 ( .B1(pipeline_md_N128), .B2(n6755), .C1(pipeline_md_N96), 
        .C2(n6754), .A(n10274), .ZN(n10281) );
  NAND2_X2 U10809 ( .A1(n6917), .A2(n10276), .ZN(n10278) );
  NOR2_X2 U10810 ( .A1(n1087), .A2(n6693), .ZN(n10279) );
  AOI221_X2 U10811 ( .B1(pipeline_md_N186), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[0]), .A(n10279), .ZN(n10280) );
  NAND2_X2 U10812 ( .A1(n10281), .A2(n10280), .ZN(n5653) );
  NAND2_X2 U10813 ( .A1(n7051), .A2(n7166), .ZN(n13115) );
  INV_X4 U10814 ( .A(n13115), .ZN(n11266) );
  NAND2_X2 U10815 ( .A1(n11229), .A2(n10282), .ZN(n10283) );
  OAI221_X2 U10816 ( .B1(n1546), .B2(n9462), .C1(n12595), .C2(n11262), .A(
        n10283), .ZN(n10284) );
  AOI221_X2 U10817 ( .B1(n11266), .B2(n10286), .C1(n11138), .C2(n10285), .A(
        n10284), .ZN(n10299) );
  OAI22_X2 U10818 ( .A1(n11264), .A2(n6828), .B1(n11269), .B2(n10287), .ZN(
        n10288) );
  AOI221_X2 U10819 ( .B1(n11136), .B2(ext_interrupts[23]), .C1(n9527), .C2(
        n10289), .A(n10288), .ZN(n10298) );
  NOR2_X2 U10820 ( .A1(n13111), .A2(n6846), .ZN(n10290) );
  AOI221_X2 U10821 ( .B1(pipeline_csr_from_host[31]), .B2(n9461), .C1(
        pipeline_csr_mscratch[31]), .C2(n11268), .A(n10290), .ZN(n10291) );
  OAI221_X2 U10822 ( .B1(n10783), .B2(n6838), .C1(n13098), .C2(n10292), .A(
        n10291), .ZN(n10296) );
  OAI22_X2 U10823 ( .A1(n9460), .A2(n10293), .B1(n9526), .B2(n6897), .ZN(
        n10295) );
  OAI22_X2 U10824 ( .A1(n13099), .A2(n6758), .B1(n13105), .B2(n6915), .ZN(
        n10294) );
  NOR3_X2 U10825 ( .A1(n10296), .A2(n10295), .A3(n10294), .ZN(n10297) );
  NOR2_X2 U10826 ( .A1(pipeline_rs1_data_bypassed[31]), .A2(n9463), .ZN(n10300) );
  NOR2_X2 U10827 ( .A1(n6793), .A2(n10300), .ZN(n10302) );
  NAND2_X2 U10828 ( .A1(htif_pcr_req_data[31]), .A2(n13131), .ZN(n10301) );
  OAI22_X2 U10829 ( .A1(n12601), .A2(n6690), .B1(n1222), .B2(n6708), .ZN(n6177) );
  OAI22_X2 U10830 ( .A1(n1546), .A2(n6660), .B1(n12601), .B2(n9516), .ZN(n6238) );
  INV_X4 U10831 ( .A(imem_hready), .ZN(n10303) );
  NAND2_X2 U10832 ( .A1(n10304), .A2(n10303), .ZN(n10305) );
  NAND3_X2 U10833 ( .A1(n10306), .A2(n13130), .A3(n10305), .ZN(
        pipeline_ctrl_N66) );
  INV_X4 U10834 ( .A(pipeline_md_N252), .ZN(n10307) );
  OAI22_X2 U10835 ( .A1(n1088), .A2(n9504), .B1(n9505), .B2(n10307), .ZN(
        n10308) );
  AOI221_X2 U10836 ( .B1(pipeline_md_N30), .B2(n6798), .C1(n6808), .C2(n6637), 
        .A(n10308), .ZN(n10309) );
  INV_X4 U10837 ( .A(n10309), .ZN(n5681) );
  INV_X4 U10838 ( .A(pipeline_md_result_muxed[33]), .ZN(n10311) );
  NOR2_X2 U10839 ( .A1(pipeline_md_N316), .A2(pipeline_md_resp_result[1]), 
        .ZN(n10310) );
  OAI22_X2 U10840 ( .A1(n10311), .A2(n6692), .B1(n10310), .B2(n6667), .ZN(
        n10312) );
  AOI221_X2 U10841 ( .B1(pipeline_md_N129), .B2(n6755), .C1(pipeline_md_N97), 
        .C2(n6754), .A(n10312), .ZN(n10315) );
  NOR2_X2 U10842 ( .A1(n1088), .A2(n6693), .ZN(n10313) );
  AOI221_X2 U10843 ( .B1(pipeline_md_N187), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[1]), .A(n10313), .ZN(n10314) );
  NAND2_X2 U10844 ( .A1(n10315), .A2(n10314), .ZN(n5652) );
  NAND2_X2 U10845 ( .A1(n10824), .A2(n13130), .ZN(n11283) );
  NAND2_X2 U10846 ( .A1(pipeline_dmem_type_2_), .A2(n6698), .ZN(n11280) );
  INV_X4 U10847 ( .A(n11280), .ZN(n10332) );
  NAND2_X2 U10848 ( .A1(pipeline_csr_time_full[33]), .A2(n11257), .ZN(n10316)
         );
  OAI221_X2 U10849 ( .B1(n13098), .B2(n10317), .C1(n13099), .C2(n6817), .A(
        n10316), .ZN(n10318) );
  AOI221_X2 U10850 ( .B1(pipeline_csr_time_full[1]), .B2(n6735), .C1(
        pipeline_csr_instret_full[1]), .C2(n6640), .A(n10318), .ZN(n10328) );
  OAI22_X2 U10851 ( .A1(n1448), .A2(n9464), .B1(n1256), .B2(n11261), .ZN(
        n10319) );
  AOI221_X2 U10852 ( .B1(pipeline_csr_from_host[1]), .B2(n9461), .C1(
        pipeline_csr_cycle_full[1]), .C2(n13116), .A(n10319), .ZN(n10327) );
  OAI22_X2 U10853 ( .A1(n11264), .A2(n6815), .B1(n1484), .B2(n13114), .ZN(
        n10320) );
  AOI221_X2 U10854 ( .B1(n11268), .B2(n10322), .C1(n11266), .C2(n10321), .A(
        n10320), .ZN(n10326) );
  NAND2_X2 U10855 ( .A1(n7063), .A2(n6641), .ZN(n13112) );
  OAI22_X2 U10856 ( .A1(n13112), .A2(n10323), .B1(n1516), .B2(n9462), .ZN(
        n10324) );
  AOI221_X2 U10857 ( .B1(pipeline_csr_mtime_full[33]), .B2(n9528), .C1(n9466), 
        .C2(pipeline_csr_mtimecmp[1]), .A(n10324), .ZN(n10325) );
  NAND4_X2 U10858 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n12391) );
  NAND2_X2 U10859 ( .A1(n6665), .A2(n12391), .ZN(n10329) );
  OAI22_X2 U10860 ( .A1(n10330), .A2(n10329), .B1(n13141), .B2(n3704), .ZN(
        n10331) );
  INV_X4 U10861 ( .A(n1911), .ZN(n12385) );
  NAND2_X2 U10862 ( .A1(n9468), .A2(n12385), .ZN(n12354) );
  NAND2_X2 U10863 ( .A1(n11318), .A2(n11282), .ZN(n10343) );
  INV_X4 U10864 ( .A(n10343), .ZN(n10335) );
  NAND4_X2 U10865 ( .A1(n7089), .A2(n10338), .A3(n9402), .A4(n10337), .ZN(
        n10350) );
  NAND3_X2 U10866 ( .A1(n7089), .A2(n6711), .A3(n9402), .ZN(n10353) );
  NAND4_X2 U10867 ( .A1(n6700), .A2(n12255), .A3(n12612), .A4(n12258), .ZN(
        n10419) );
  NAND2_X2 U10868 ( .A1(n6714), .A2(n6749), .ZN(n10340) );
  NAND2_X2 U10869 ( .A1(n9468), .A2(n10340), .ZN(n10342) );
  NAND2_X2 U10870 ( .A1(n10341), .A2(n13130), .ZN(n11320) );
  NAND2_X2 U10871 ( .A1(n10342), .A2(n11320), .ZN(n11198) );
  INV_X4 U10872 ( .A(pipeline_csr_N745), .ZN(n10344) );
  OAI22_X2 U10873 ( .A1(n9492), .A2(n12354), .B1(n9403), .B2(n10344), .ZN(
        pipeline_csr_N1985) );
  NAND2_X2 U10874 ( .A1(n12395), .A2(n13130), .ZN(n11179) );
  NOR2_X2 U10875 ( .A1(pipeline_ctrl_prev_killed_DX), .A2(n10346), .ZN(n10347)
         );
  OAI22_X2 U10876 ( .A1(n10347), .A2(n12827), .B1(n793), .B2(n12829), .ZN(
        n6048) );
  INV_X4 U10877 ( .A(n10350), .ZN(n10522) );
  NAND2_X2 U10878 ( .A1(n10522), .A2(n10824), .ZN(n10351) );
  NAND2_X2 U10879 ( .A1(n9468), .A2(n12352), .ZN(n10354) );
  INV_X4 U10880 ( .A(n10354), .ZN(n10352) );
  INV_X4 U10881 ( .A(n10353), .ZN(n10519) );
  NAND2_X2 U10882 ( .A1(n6714), .A2(n6820), .ZN(n10521) );
  NOR2_X2 U10883 ( .A1(n10519), .A2(n10521), .ZN(n10355) );
  OAI22_X2 U10884 ( .A1(n10355), .A2(n10354), .B1(n9478), .B2(n11320), .ZN(
        n12350) );
  NAND2_X2 U10885 ( .A1(pipeline_csr_N839), .A2(n9476), .ZN(n10356) );
  OAI221_X2 U10886 ( .B1(n12601), .B2(n6704), .C1(n10292), .C2(n12352), .A(
        n10356), .ZN(n5984) );
  NAND2_X2 U10887 ( .A1(pipeline_csr_N838), .A2(n9476), .ZN(n10357) );
  OAI221_X2 U10888 ( .B1(n12670), .B2(n6704), .C1(n1445), .C2(n12352), .A(
        n10357), .ZN(n5985) );
  NAND2_X2 U10889 ( .A1(n11229), .A2(n10358), .ZN(n10359) );
  OAI221_X2 U10890 ( .B1(n1544), .B2(n9462), .C1(n12328), .C2(n11262), .A(
        n10359), .ZN(n10360) );
  AOI221_X2 U10891 ( .B1(n11138), .B2(n10361), .C1(n11136), .C2(
        ext_interrupts[21]), .A(n10360), .ZN(n10372) );
  OAI22_X2 U10892 ( .A1(n13111), .A2(n6867), .B1(n11269), .B2(n10362), .ZN(
        n10363) );
  AOI221_X2 U10893 ( .B1(n9527), .B2(n10364), .C1(pipeline_csr_mtime_full[29]), 
        .C2(n13108), .A(n10363), .ZN(n10371) );
  OAI22_X2 U10894 ( .A1(n13105), .A2(n6868), .B1(n11235), .B2(n10365), .ZN(
        n10366) );
  AOI221_X2 U10895 ( .B1(pipeline_csr_mscratch[29]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[29]), .C2(n13116), .A(n10366), .ZN(n10370) );
  OAI22_X2 U10896 ( .A1(n9526), .A2(n6887), .B1(n9460), .B2(n10367), .ZN(
        n10368) );
  AOI221_X2 U10897 ( .B1(pipeline_csr_instret_full[61]), .B2(n11105), .C1(
        pipeline_csr_cycle_full[61]), .C2(n11233), .A(n10368), .ZN(n10369) );
  NOR2_X2 U10898 ( .A1(pipeline_rs1_data_bypassed[29]), .A2(n9463), .ZN(n10373) );
  NOR2_X2 U10899 ( .A1(n6793), .A2(n10373), .ZN(n10375) );
  NAND2_X2 U10900 ( .A1(htif_pcr_req_data[29]), .A2(n13131), .ZN(n10374) );
  OAI221_X2 U10901 ( .B1(n7210), .B2(n10375), .C1(n12422), .C2(n9467), .A(
        n10374), .ZN(n12330) );
  INV_X4 U10902 ( .A(n12330), .ZN(n12338) );
  OAI22_X2 U10903 ( .A1(n12338), .A2(n6690), .B1(n1220), .B2(n6708), .ZN(n6179) );
  OAI22_X2 U10904 ( .A1(n12338), .A2(n9516), .B1(n1544), .B2(n6660), .ZN(n6236) );
  INV_X4 U10905 ( .A(pipeline_md_N280), .ZN(n10376) );
  OAI22_X2 U10906 ( .A1(n1116), .A2(n9504), .B1(n12765), .B2(n10376), .ZN(
        n10377) );
  INV_X4 U10907 ( .A(n10378), .ZN(n5682) );
  INV_X4 U10908 ( .A(pipeline_md_result_muxed[61]), .ZN(n10380) );
  NOR2_X2 U10909 ( .A1(pipeline_md_N344), .A2(pipeline_md_resp_result[29]), 
        .ZN(n10379) );
  OAI22_X2 U10910 ( .A1(n10380), .A2(n6692), .B1(n10379), .B2(n6667), .ZN(
        n10381) );
  AOI221_X2 U10911 ( .B1(pipeline_md_N157), .B2(n6755), .C1(pipeline_md_N125), 
        .C2(n6754), .A(n10381), .ZN(n10384) );
  NOR2_X2 U10912 ( .A1(n1116), .A2(n6693), .ZN(n10382) );
  AOI221_X2 U10913 ( .B1(pipeline_md_N215), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[29]), .A(n10382), .ZN(n10383) );
  NAND2_X2 U10914 ( .A1(n10384), .A2(n10383), .ZN(n5624) );
  OAI22_X2 U10915 ( .A1(n7210), .A2(n6691), .B1(n466), .B2(n9523), .ZN(n6363)
         );
  INV_X4 U10916 ( .A(n10385), .ZN(n10386) );
  NAND2_X2 U10917 ( .A1(n9493), .A2(n13130), .ZN(n12632) );
  INV_X4 U10918 ( .A(n13162), .ZN(n10387) );
  OAI22_X2 U10919 ( .A1(n12425), .A2(n9494), .B1(n9493), .B2(n10387), .ZN(
        n5942) );
  OAI22_X2 U10920 ( .A1(n12425), .A2(n9496), .B1(n744), .B2(n6662), .ZN(n5881)
         );
  INV_X4 U10921 ( .A(pipeline_md_N253), .ZN(n10389) );
  OAI22_X2 U10922 ( .A1(n13046), .A2(n9504), .B1(n9505), .B2(n10389), .ZN(
        n10390) );
  INV_X4 U10923 ( .A(n10391), .ZN(n5654) );
  INV_X4 U10924 ( .A(pipeline_md_result_muxed[34]), .ZN(n10393) );
  NOR2_X2 U10925 ( .A1(pipeline_md_N317), .A2(pipeline_md_resp_result[2]), 
        .ZN(n10392) );
  OAI22_X2 U10926 ( .A1(n10393), .A2(n6692), .B1(n10392), .B2(n6667), .ZN(
        n10394) );
  AOI221_X2 U10927 ( .B1(pipeline_md_N130), .B2(n6755), .C1(pipeline_md_N98), 
        .C2(n6754), .A(n10394), .ZN(n10397) );
  NOR2_X2 U10928 ( .A1(n13046), .A2(n6693), .ZN(n10395) );
  AOI221_X2 U10929 ( .B1(pipeline_md_N188), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[2]), .A(n10395), .ZN(n10396) );
  NAND2_X2 U10930 ( .A1(n10397), .A2(n10396), .ZN(n5651) );
  NAND2_X2 U10931 ( .A1(pipeline_csr_mtvec[2]), .A2(n11229), .ZN(n10398) );
  OAI221_X2 U10932 ( .B1(n13105), .B2(n6835), .C1(n13098), .C2(n10399), .A(
        n10398), .ZN(n10400) );
  AOI221_X2 U10933 ( .B1(pipeline_csr_cycle_full[34]), .B2(n11233), .C1(
        pipeline_csr_time_full[2]), .C2(n6735), .A(n10400), .ZN(n10412) );
  OAI22_X2 U10934 ( .A1(n11235), .A2(n10401), .B1(n12288), .B2(n9464), .ZN(
        n10402) );
  AOI221_X2 U10935 ( .B1(pipeline_csr_instret_full[2]), .B2(n6640), .C1(n9527), 
        .C2(n10403), .A(n10402), .ZN(n10411) );
  NAND2_X2 U10936 ( .A1(pipeline_csr_cycle_full[2]), .A2(n13116), .ZN(n10404)
         );
  OAI221_X2 U10937 ( .B1(n1163), .B2(n13113), .C1(n1481), .C2(n13115), .A(
        n10404), .ZN(n10405) );
  AOI221_X2 U10938 ( .B1(n11138), .B2(n10406), .C1(pipeline_csr_mtime_full[2]), 
        .C2(n13108), .A(n10405), .ZN(n10410) );
  OAI22_X2 U10939 ( .A1(n13112), .A2(n10407), .B1(n1517), .B2(n9462), .ZN(
        n10408) );
  AOI221_X2 U10940 ( .B1(pipeline_csr_mtime_full[34]), .B2(n9528), .C1(n9466), 
        .C2(pipeline_csr_mtimecmp[2]), .A(n10408), .ZN(n10409) );
  NAND4_X2 U10941 ( .A1(n10412), .A2(n10411), .A3(n10410), .A4(n10409), .ZN(
        n12295) );
  NAND2_X2 U10942 ( .A1(n6665), .A2(n12295), .ZN(n10413) );
  OAI22_X2 U10943 ( .A1(n1909), .A2(n6690), .B1(n1193), .B2(n6708), .ZN(n6206)
         );
  NAND2_X2 U10944 ( .A1(n9468), .A2(n10416), .ZN(n12260) );
  INV_X4 U10945 ( .A(pipeline_csr_N746), .ZN(n10417) );
  OAI22_X2 U10946 ( .A1(n9492), .A2(n12260), .B1(n9403), .B2(n10417), .ZN(
        pipeline_csr_N1986) );
  NAND2_X2 U10947 ( .A1(pipeline_csr_N810), .A2(n9476), .ZN(n10418) );
  OAI221_X2 U10948 ( .B1(n1909), .B2(n6704), .C1(n10399), .C2(n12352), .A(
        n10418), .ZN(n6012) );
  NAND3_X2 U10949 ( .A1(n10419), .A2(n12255), .A3(n6700), .ZN(n10420) );
  NAND2_X2 U10950 ( .A1(n9468), .A2(n10420), .ZN(n10421) );
  NAND2_X2 U10951 ( .A1(n10421), .A2(n11320), .ZN(n10516) );
  INV_X4 U10952 ( .A(pipeline_csr_N711), .ZN(n10423) );
  NAND2_X2 U10953 ( .A1(n9468), .A2(n10422), .ZN(n12603) );
  OAI22_X2 U10954 ( .A1(n12257), .A2(n10423), .B1(n9469), .B2(n12603), .ZN(
        pipeline_csr_N1951) );
  NAND2_X2 U10955 ( .A1(n9468), .A2(n12667), .ZN(n12607) );
  INV_X4 U10956 ( .A(pipeline_csr_N710), .ZN(n10424) );
  OAI22_X2 U10957 ( .A1(n9469), .A2(n12607), .B1(n9404), .B2(n10424), .ZN(
        pipeline_csr_N1950) );
  NAND2_X2 U10958 ( .A1(n9468), .A2(n12330), .ZN(n12335) );
  INV_X4 U10959 ( .A(pipeline_csr_N709), .ZN(n10425) );
  OAI22_X2 U10960 ( .A1(n9469), .A2(n12335), .B1(n12257), .B2(n10425), .ZN(
        pipeline_csr_N1949) );
  NAND2_X2 U10961 ( .A1(n11229), .A2(n10426), .ZN(n10427) );
  OAI221_X2 U10962 ( .B1(n1543), .B2(n9462), .C1(n12232), .C2(n11262), .A(
        n10427), .ZN(n10428) );
  AOI221_X2 U10963 ( .B1(n11138), .B2(n10429), .C1(n11136), .C2(
        ext_interrupts[20]), .A(n10428), .ZN(n10438) );
  OAI22_X2 U10964 ( .A1(n11269), .A2(n10430), .B1(n1283), .B2(n11261), .ZN(
        n10431) );
  AOI221_X2 U10965 ( .B1(pipeline_csr_mtime_full[28]), .B2(n13108), .C1(
        pipeline_csr_mscratch[28]), .C2(n11268), .A(n10431), .ZN(n10437) );
  OAI22_X2 U10966 ( .A1(n13099), .A2(n6869), .B1(n10783), .B2(n6752), .ZN(
        n10432) );
  OAI22_X2 U10967 ( .A1(n9460), .A2(n10433), .B1(n9526), .B2(n6831), .ZN(
        n10434) );
  AOI221_X2 U10968 ( .B1(pipeline_csr_time_full[60]), .B2(n11257), .C1(
        pipeline_csr_instret_full[60]), .C2(n11105), .A(n10434), .ZN(n10435)
         );
  NOR2_X2 U10969 ( .A1(pipeline_rs1_data_bypassed[28]), .A2(n9463), .ZN(n10439) );
  NOR2_X2 U10970 ( .A1(n6793), .A2(n10439), .ZN(n10441) );
  NAND2_X2 U10971 ( .A1(htif_pcr_req_data[28]), .A2(n13131), .ZN(n10440) );
  OAI221_X2 U10972 ( .B1(n7212), .B2(n10441), .C1(n12426), .C2(n9467), .A(
        n10440), .ZN(n12234) );
  INV_X4 U10973 ( .A(n12234), .ZN(n12242) );
  OAI22_X2 U10974 ( .A1(n12242), .A2(n6690), .B1(n1219), .B2(n6708), .ZN(n6180) );
  OAI22_X2 U10975 ( .A1(n12242), .A2(n9516), .B1(n1543), .B2(n6660), .ZN(n6235) );
  INV_X4 U10976 ( .A(pipeline_md_N279), .ZN(n10442) );
  AOI221_X2 U10978 ( .B1(pipeline_md_N57), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[28]), .A(n10443), .ZN(n10444) );
  INV_X4 U10979 ( .A(n10444), .ZN(n5680) );
  INV_X4 U10980 ( .A(pipeline_md_result_muxed[60]), .ZN(n10446) );
  NOR2_X2 U10981 ( .A1(pipeline_md_N343), .A2(pipeline_md_resp_result[28]), 
        .ZN(n10445) );
  OAI22_X2 U10982 ( .A1(n10446), .A2(n6692), .B1(n10445), .B2(n6667), .ZN(
        n10447) );
  AOI221_X2 U10983 ( .B1(pipeline_md_N156), .B2(n6755), .C1(pipeline_md_N124), 
        .C2(n6754), .A(n10447), .ZN(n10450) );
  NOR2_X2 U10984 ( .A1(n1115), .A2(n6693), .ZN(n10448) );
  AOI221_X2 U10985 ( .B1(pipeline_md_N214), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[28]), .A(n10448), .ZN(n10449) );
  NAND2_X2 U10986 ( .A1(n10450), .A2(n10449), .ZN(n5625) );
  OAI22_X2 U10987 ( .A1(n7212), .A2(n6691), .B1(n464), .B2(n9524), .ZN(n6362)
         );
  INV_X4 U10988 ( .A(n13163), .ZN(n10451) );
  OAI22_X2 U10989 ( .A1(n12429), .A2(n12632), .B1(n9493), .B2(n10451), .ZN(
        n5943) );
  OAI22_X2 U10990 ( .A1(n12429), .A2(n9496), .B1(n743), .B2(n6662), .ZN(n5883)
         );
  INV_X4 U10991 ( .A(pipeline_md_N278), .ZN(n10452) );
  OAI22_X2 U10992 ( .A1(n13054), .A2(n9504), .B1(n12765), .B2(n10452), .ZN(
        n10453) );
  INV_X4 U10993 ( .A(n10454), .ZN(n5679) );
  INV_X4 U10994 ( .A(pipeline_md_result_muxed[59]), .ZN(n10456) );
  NOR2_X2 U10995 ( .A1(pipeline_md_N342), .A2(pipeline_md_resp_result[27]), 
        .ZN(n10455) );
  OAI22_X2 U10996 ( .A1(n10456), .A2(n6692), .B1(n10455), .B2(n6667), .ZN(
        n10457) );
  AOI221_X2 U10997 ( .B1(pipeline_md_N155), .B2(n6755), .C1(pipeline_md_N123), 
        .C2(n6754), .A(n10457), .ZN(n10460) );
  NOR2_X2 U10998 ( .A1(n13054), .A2(n6693), .ZN(n10458) );
  AOI221_X2 U10999 ( .B1(pipeline_md_N213), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[27]), .A(n10458), .ZN(n10459) );
  NAND2_X2 U11000 ( .A1(n10460), .A2(n10459), .ZN(n5626) );
  NAND2_X2 U11001 ( .A1(n11229), .A2(n10461), .ZN(n10462) );
  OAI221_X2 U11002 ( .B1(n1542), .B2(n9462), .C1(n12186), .C2(n11262), .A(
        n10462), .ZN(n10463) );
  AOI221_X2 U11003 ( .B1(n11138), .B2(n10464), .C1(n11136), .C2(
        ext_interrupts[19]), .A(n10463), .ZN(n10475) );
  OAI22_X2 U11004 ( .A1(n13111), .A2(n6870), .B1(n11269), .B2(n10465), .ZN(
        n10466) );
  AOI221_X2 U11005 ( .B1(n9527), .B2(n10467), .C1(pipeline_csr_mtime_full[27]), 
        .C2(n13108), .A(n10466), .ZN(n10474) );
  OAI22_X2 U11006 ( .A1(n13105), .A2(n6871), .B1(n11235), .B2(n10468), .ZN(
        n10469) );
  AOI221_X2 U11007 ( .B1(pipeline_csr_mscratch[27]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[27]), .C2(n13116), .A(n10469), .ZN(n10473) );
  OAI22_X2 U11008 ( .A1(n9460), .A2(n10470), .B1(n9526), .B2(n6898), .ZN(
        n10471) );
  AOI221_X2 U11009 ( .B1(pipeline_csr_cycle_full[59]), .B2(n11233), .C1(
        pipeline_csr_instret_full[59]), .C2(n11105), .A(n10471), .ZN(n10472)
         );
  NOR2_X2 U11010 ( .A1(n6793), .A2(n10476), .ZN(n10478) );
  NAND2_X2 U11011 ( .A1(htif_pcr_req_data[27]), .A2(n13131), .ZN(n10477) );
  OAI221_X2 U11012 ( .B1(n7209), .B2(n10478), .C1(n12430), .C2(n9467), .A(
        n10477), .ZN(n12188) );
  INV_X4 U11013 ( .A(n12188), .ZN(n12198) );
  OAI22_X2 U11014 ( .A1(n12198), .A2(n6690), .B1(n1218), .B2(n6708), .ZN(n6181) );
  OAI22_X2 U11015 ( .A1(n12198), .A2(n9516), .B1(n1542), .B2(n6660), .ZN(n6234) );
  INV_X4 U11016 ( .A(pipeline_md_N254), .ZN(n10479) );
  OAI22_X2 U11017 ( .A1(n13045), .A2(n9504), .B1(n9505), .B2(n10479), .ZN(
        n10480) );
  INV_X4 U11018 ( .A(n10481), .ZN(n5655) );
  INV_X4 U11019 ( .A(pipeline_md_result_muxed[35]), .ZN(n10483) );
  NOR2_X2 U11020 ( .A1(pipeline_md_N318), .A2(pipeline_md_resp_result[3]), 
        .ZN(n10482) );
  OAI22_X2 U11021 ( .A1(n10483), .A2(n6692), .B1(n10482), .B2(n6667), .ZN(
        n10484) );
  AOI221_X2 U11022 ( .B1(pipeline_md_N131), .B2(n6755), .C1(pipeline_md_N99), 
        .C2(n6754), .A(n10484), .ZN(n10487) );
  NOR2_X2 U11023 ( .A1(n13045), .A2(n6693), .ZN(n10485) );
  AOI221_X2 U11024 ( .B1(pipeline_md_N189), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[3]), .A(n10485), .ZN(n10486) );
  NAND2_X2 U11025 ( .A1(n10487), .A2(n10486), .ZN(n5650) );
  NAND2_X2 U11026 ( .A1(htif_pcr_req_data[3]), .A2(n13131), .ZN(n10509) );
  NAND2_X2 U11027 ( .A1(pipeline_regfile_N15), .A2(pipeline_dmem_type_2_), 
        .ZN(n10504) );
  NAND2_X2 U11028 ( .A1(n11136), .A2(pipeline_csr_mip_3), .ZN(n10488) );
  OAI221_X2 U11029 ( .B1(n13104), .B2(n10489), .C1(n13105), .C2(n6837), .A(
        n10488), .ZN(n10490) );
  AOI221_X2 U11030 ( .B1(pipeline_csr_instret_full[35]), .B2(n11105), .C1(
        pipeline_csr_cycle_full[35]), .C2(n11233), .A(n10490), .ZN(n10501) );
  NAND2_X2 U11031 ( .A1(pipeline_csr_to_host_3_), .A2(n9527), .ZN(n10491) );
  OAI221_X2 U11032 ( .B1(n9526), .B2(n6839), .C1(n9460), .C2(n10492), .A(
        n10491), .ZN(n10493) );
  AOI221_X2 U11033 ( .B1(pipeline_csr_mbadaddr[3]), .B2(n9465), .C1(
        pipeline_csr_from_host[3]), .C2(n9461), .A(n10493), .ZN(n10500) );
  NAND2_X2 U11034 ( .A1(pipeline_csr_cycle_full[3]), .A2(n13116), .ZN(n10494)
         );
  OAI221_X2 U11035 ( .B1(n1164), .B2(n13113), .C1(n1482), .C2(n13115), .A(
        n10494), .ZN(n10495) );
  AOI221_X2 U11036 ( .B1(n11138), .B2(n10496), .C1(pipeline_csr_mtime_full[3]), 
        .C2(n13108), .A(n10495), .ZN(n10499) );
  OAI22_X2 U11037 ( .A1(n13112), .A2(n12155), .B1(n1518), .B2(n9462), .ZN(
        n10497) );
  AOI221_X2 U11038 ( .B1(pipeline_csr_mtime_full[35]), .B2(n9528), .C1(n9466), 
        .C2(pipeline_csr_mtimecmp[3]), .A(n10497), .ZN(n10498) );
  NOR2_X2 U11039 ( .A1(n6701), .A2(n9463), .ZN(n10503) );
  NAND3_X2 U11040 ( .A1(n10504), .A2(n10503), .A3(n10502), .ZN(n10508) );
  NOR2_X2 U11041 ( .A1(n12526), .A2(n9467), .ZN(n10506) );
  NOR2_X2 U11042 ( .A1(n11280), .A2(n9279), .ZN(n10505) );
  NOR2_X2 U11043 ( .A1(n10506), .A2(n10505), .ZN(n10507) );
  NAND3_X2 U11044 ( .A1(n10509), .A2(n10508), .A3(n10507), .ZN(n10512) );
  INV_X4 U11045 ( .A(n10512), .ZN(n1907) );
  MUX2_X2 U11046 ( .A(n10510), .B(n1907), .S(n6826), .Z(n10511) );
  NOR2_X2 U11047 ( .A1(htif_reset), .A2(n10511), .ZN(n6240) );
  OAI22_X2 U11048 ( .A1(n1907), .A2(n6690), .B1(n10489), .B2(n6708), .ZN(n6205) );
  NAND2_X2 U11049 ( .A1(n9468), .A2(n10512), .ZN(n12147) );
  INV_X4 U11050 ( .A(pipeline_csr_N747), .ZN(n10513) );
  OAI22_X2 U11051 ( .A1(n9492), .A2(n12147), .B1(n9403), .B2(n10513), .ZN(
        pipeline_csr_N1987) );
  NAND2_X2 U11052 ( .A1(pipeline_csr_N811), .A2(n9476), .ZN(n10514) );
  OAI221_X2 U11053 ( .B1(n1907), .B2(n6704), .C1(n1418), .C2(n12352), .A(
        n10514), .ZN(n6011) );
  INV_X4 U11054 ( .A(pipeline_csr_N683), .ZN(n10515) );
  OAI22_X2 U11055 ( .A1(n9469), .A2(n12147), .B1(n12257), .B2(n10515), .ZN(
        pipeline_csr_N1923) );
  INV_X4 U11056 ( .A(pipeline_csr_N715), .ZN(n10517) );
  OAI22_X2 U11057 ( .A1(n12612), .A2(n12147), .B1(n9405), .B2(n10517), .ZN(
        pipeline_csr_N1955) );
  NAND2_X2 U11058 ( .A1(n10519), .A2(n10824), .ZN(n10518) );
  NAND2_X2 U11059 ( .A1(n9468), .A2(n12349), .ZN(n10523) );
  INV_X4 U11060 ( .A(n10523), .ZN(n10520) );
  NOR2_X2 U11061 ( .A1(n10522), .A2(n10521), .ZN(n10524) );
  OAI22_X2 U11062 ( .A1(n10524), .A2(n10523), .B1(n9475), .B2(n11320), .ZN(
        n12346) );
  NAND2_X2 U11063 ( .A1(pipeline_csr_N779), .A2(n9472), .ZN(n10525) );
  OAI221_X2 U11064 ( .B1(n1907), .B2(n12347), .C1(n10492), .C2(n12349), .A(
        n10525), .ZN(n6043) );
  INV_X4 U11065 ( .A(imem_haddr[3]), .ZN(n10526) );
  OAI22_X2 U11066 ( .A1(n12529), .A2(n12632), .B1(n9493), .B2(n10526), .ZN(
        n5968) );
  OAI22_X2 U11067 ( .A1(n12529), .A2(n9496), .B1(n718), .B2(n6662), .ZN(n5933)
         );
  INV_X4 U11068 ( .A(imem_haddr[2]), .ZN(n10527) );
  OAI22_X2 U11069 ( .A1(n12534), .A2(n12632), .B1(n9493), .B2(n10527), .ZN(
        n5969) );
  OAI22_X2 U11070 ( .A1(n12534), .A2(n9496), .B1(n717), .B2(n6662), .ZN(n5935)
         );
  INV_X4 U11071 ( .A(pipeline_md_N277), .ZN(n10528) );
  AOI221_X2 U11073 ( .B1(pipeline_md_N55), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[26]), .A(n10529), .ZN(n10530) );
  INV_X4 U11074 ( .A(n10530), .ZN(n5678) );
  INV_X4 U11075 ( .A(pipeline_md_result_muxed[58]), .ZN(n10532) );
  NOR2_X2 U11076 ( .A1(pipeline_md_N341), .A2(pipeline_md_resp_result[26]), 
        .ZN(n10531) );
  OAI22_X2 U11077 ( .A1(n10532), .A2(n6692), .B1(n10531), .B2(n6667), .ZN(
        n10533) );
  AOI221_X2 U11078 ( .B1(pipeline_md_N154), .B2(n6755), .C1(pipeline_md_N122), 
        .C2(n6754), .A(n10533), .ZN(n10536) );
  NOR2_X2 U11079 ( .A1(n13055), .A2(n6693), .ZN(n10534) );
  AOI221_X2 U11080 ( .B1(pipeline_md_N212), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[26]), .A(n10534), .ZN(n10535) );
  NAND2_X2 U11081 ( .A1(n10536), .A2(n10535), .ZN(n5627) );
  NAND2_X2 U11082 ( .A1(n11229), .A2(n10537), .ZN(n10538) );
  OAI221_X2 U11083 ( .B1(n1541), .B2(n9462), .C1(n12108), .C2(n9464), .A(
        n10538), .ZN(n10539) );
  AOI221_X2 U11084 ( .B1(n11138), .B2(n10540), .C1(n11136), .C2(
        ext_interrupts[18]), .A(n10539), .ZN(n10551) );
  OAI22_X2 U11085 ( .A1(n13111), .A2(n6872), .B1(n11269), .B2(n10541), .ZN(
        n10542) );
  AOI221_X2 U11086 ( .B1(n9527), .B2(n10543), .C1(pipeline_csr_mtime_full[26]), 
        .C2(n13108), .A(n10542), .ZN(n10550) );
  OAI22_X2 U11087 ( .A1(n13105), .A2(n6873), .B1(n11235), .B2(n10544), .ZN(
        n10545) );
  AOI221_X2 U11088 ( .B1(pipeline_csr_mscratch[26]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[26]), .C2(n13116), .A(n10545), .ZN(n10549) );
  OAI22_X2 U11089 ( .A1(n9460), .A2(n10546), .B1(n9526), .B2(n6832), .ZN(
        n10547) );
  AOI221_X2 U11090 ( .B1(pipeline_csr_cycle_full[58]), .B2(n11233), .C1(
        pipeline_csr_instret_full[58]), .C2(n11105), .A(n10547), .ZN(n10548)
         );
  NOR2_X2 U11091 ( .A1(pipeline_rs1_data_bypassed[26]), .A2(n9463), .ZN(n10552) );
  NOR2_X2 U11092 ( .A1(n6793), .A2(n10552), .ZN(n10554) );
  NAND2_X2 U11093 ( .A1(htif_pcr_req_data[26]), .A2(n13131), .ZN(n10553) );
  OAI221_X2 U11094 ( .B1(n7208), .B2(n10554), .C1(n12434), .C2(n9467), .A(
        n10553), .ZN(n12110) );
  INV_X4 U11095 ( .A(n12110), .ZN(n12120) );
  OAI22_X2 U11096 ( .A1(n12120), .A2(n6690), .B1(n1217), .B2(n6708), .ZN(n6182) );
  OAI22_X2 U11097 ( .A1(n12120), .A2(n9516), .B1(n1541), .B2(n6660), .ZN(n6233) );
  INV_X4 U11098 ( .A(pipeline_md_N260), .ZN(n10555) );
  OAI22_X2 U11099 ( .A1(n1096), .A2(n9504), .B1(n12765), .B2(n10555), .ZN(
        n10556) );
  INV_X4 U11100 ( .A(n10557), .ZN(n5661) );
  INV_X4 U11101 ( .A(pipeline_md_result_muxed[41]), .ZN(n10559) );
  NOR2_X2 U11102 ( .A1(pipeline_md_N324), .A2(pipeline_md_resp_result[9]), 
        .ZN(n10558) );
  OAI22_X2 U11103 ( .A1(n10559), .A2(n6692), .B1(n10558), .B2(n6667), .ZN(
        n10560) );
  AOI221_X2 U11104 ( .B1(pipeline_md_N137), .B2(n6755), .C1(pipeline_md_N105), 
        .C2(n6754), .A(n10560), .ZN(n10563) );
  NOR2_X2 U11105 ( .A1(n1096), .A2(n6693), .ZN(n10561) );
  AOI221_X2 U11106 ( .B1(pipeline_md_N195), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[9]), .A(n10561), .ZN(n10562) );
  NAND2_X2 U11107 ( .A1(n10563), .A2(n10562), .ZN(n5644) );
  NAND2_X2 U11108 ( .A1(n11229), .A2(n10564), .ZN(n10565) );
  OAI221_X2 U11109 ( .B1(n1524), .B2(n9462), .C1(n12072), .C2(n11262), .A(
        n10565), .ZN(n10566) );
  AOI221_X2 U11110 ( .B1(n11138), .B2(n10567), .C1(n11136), .C2(
        ext_interrupts[1]), .A(n10566), .ZN(n10579) );
  OAI22_X2 U11111 ( .A1(n13111), .A2(n6888), .B1(n11269), .B2(n10568), .ZN(
        n10569) );
  AOI221_X2 U11112 ( .B1(n9527), .B2(n10570), .C1(pipeline_csr_mtime_full[9]), 
        .C2(n13108), .A(n10569), .ZN(n10578) );
  OAI22_X2 U11113 ( .A1(n13098), .A2(n10572), .B1(n11235), .B2(n10571), .ZN(
        n10573) );
  AOI221_X2 U11114 ( .B1(pipeline_csr_mscratch[9]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[9]), .C2(n13116), .A(n10573), .ZN(n10577) );
  OAI22_X2 U11115 ( .A1(n9526), .A2(n6889), .B1(n9460), .B2(n10574), .ZN(
        n10575) );
  AOI221_X2 U11116 ( .B1(pipeline_csr_time_full[41]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[41]), .C2(n11233), .A(n10575), .ZN(n10576) );
  NOR2_X2 U11117 ( .A1(n6793), .A2(n10580), .ZN(n10581) );
  OAI221_X2 U11118 ( .B1(n7202), .B2(n10581), .C1(n12501), .C2(n9467), .A(
        n3721), .ZN(n12074) );
  INV_X4 U11119 ( .A(n12074), .ZN(n12082) );
  OAI22_X2 U11120 ( .A1(n12082), .A2(n6690), .B1(n1200), .B2(n6708), .ZN(n6199) );
  OAI22_X2 U11121 ( .A1(n12082), .A2(n9516), .B1(n1524), .B2(n6660), .ZN(n6216) );
  INV_X4 U11122 ( .A(pipeline_md_N276), .ZN(n10582) );
  OAI22_X2 U11123 ( .A1(n1112), .A2(n9504), .B1(n12765), .B2(n10582), .ZN(
        n10583) );
  AOI221_X2 U11124 ( .B1(pipeline_md_N54), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[25]), .A(n10583), .ZN(n10584) );
  INV_X4 U11125 ( .A(n10584), .ZN(n5677) );
  INV_X4 U11126 ( .A(pipeline_md_result_muxed[57]), .ZN(n10586) );
  NOR2_X2 U11127 ( .A1(pipeline_md_N340), .A2(pipeline_md_resp_result[25]), 
        .ZN(n10585) );
  OAI22_X2 U11128 ( .A1(n10586), .A2(n6692), .B1(n10585), .B2(n6667), .ZN(
        n10587) );
  AOI221_X2 U11129 ( .B1(pipeline_md_N153), .B2(n6755), .C1(pipeline_md_N121), 
        .C2(n6754), .A(n10587), .ZN(n10590) );
  NOR2_X2 U11130 ( .A1(n1112), .A2(n6693), .ZN(n10588) );
  AOI221_X2 U11131 ( .B1(pipeline_md_N211), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[25]), .A(n10588), .ZN(n10589) );
  NAND2_X2 U11132 ( .A1(n10590), .A2(n10589), .ZN(n5628) );
  NAND2_X2 U11133 ( .A1(n11229), .A2(n10591), .ZN(n10592) );
  OAI221_X2 U11134 ( .B1(n1540), .B2(n9462), .C1(n12040), .C2(n9464), .A(
        n10592), .ZN(n10593) );
  AOI221_X2 U11135 ( .B1(n11138), .B2(n10594), .C1(n11136), .C2(
        ext_interrupts[17]), .A(n10593), .ZN(n10605) );
  OAI22_X2 U11136 ( .A1(n13111), .A2(n6874), .B1(n11269), .B2(n10595), .ZN(
        n10596) );
  AOI221_X2 U11137 ( .B1(n9527), .B2(n10597), .C1(pipeline_csr_mtime_full[25]), 
        .C2(n13108), .A(n10596), .ZN(n10604) );
  OAI22_X2 U11138 ( .A1(n13105), .A2(n6875), .B1(n11235), .B2(n10598), .ZN(
        n10599) );
  AOI221_X2 U11139 ( .B1(pipeline_csr_mscratch[25]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[25]), .C2(n13116), .A(n10599), .ZN(n10603) );
  OAI22_X2 U11140 ( .A1(n9460), .A2(n10600), .B1(n9526), .B2(n6899), .ZN(
        n10601) );
  AOI221_X2 U11141 ( .B1(pipeline_csr_cycle_full[57]), .B2(n11233), .C1(
        pipeline_csr_instret_full[57]), .C2(n11105), .A(n10601), .ZN(n10602)
         );
  NOR2_X2 U11142 ( .A1(pipeline_rs1_data_bypassed[25]), .A2(n9463), .ZN(n10606) );
  NOR2_X2 U11143 ( .A1(n6793), .A2(n10606), .ZN(n10608) );
  NAND2_X2 U11144 ( .A1(htif_pcr_req_data[25]), .A2(n13131), .ZN(n10607) );
  OAI221_X2 U11145 ( .B1(n7207), .B2(n10608), .C1(n12438), .C2(n9467), .A(
        n10607), .ZN(n12042) );
  INV_X4 U11146 ( .A(n12042), .ZN(n12052) );
  OAI22_X2 U11147 ( .A1(n12052), .A2(n6690), .B1(n1216), .B2(n6708), .ZN(n6183) );
  OAI22_X2 U11148 ( .A1(n12052), .A2(n9516), .B1(n1540), .B2(n6660), .ZN(n6232) );
  INV_X4 U11149 ( .A(pipeline_md_N259), .ZN(n10609) );
  OAI22_X2 U11150 ( .A1(n1095), .A2(n9504), .B1(n12765), .B2(n10609), .ZN(
        n10610) );
  INV_X4 U11151 ( .A(n10611), .ZN(n5660) );
  INV_X4 U11152 ( .A(pipeline_md_result_muxed[40]), .ZN(n10613) );
  NOR2_X2 U11153 ( .A1(pipeline_md_N323), .A2(pipeline_md_resp_result[8]), 
        .ZN(n10612) );
  OAI22_X2 U11154 ( .A1(n10613), .A2(n6692), .B1(n10612), .B2(n6667), .ZN(
        n10614) );
  AOI221_X2 U11155 ( .B1(pipeline_md_N136), .B2(n6755), .C1(pipeline_md_N104), 
        .C2(n6754), .A(n10614), .ZN(n10617) );
  NOR2_X2 U11156 ( .A1(n1095), .A2(n6693), .ZN(n10615) );
  AOI221_X2 U11157 ( .B1(pipeline_md_N194), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[8]), .A(n10615), .ZN(n10616) );
  NAND2_X2 U11158 ( .A1(n10617), .A2(n10616), .ZN(n5645) );
  NAND2_X2 U11159 ( .A1(n11105), .A2(n10618), .ZN(n10619) );
  OAI221_X2 U11160 ( .B1(n11264), .B2(n6825), .C1(n11269), .C2(n10620), .A(
        n10619), .ZN(n10621) );
  AOI221_X2 U11161 ( .B1(pipeline_csr_mtime_full[40]), .B2(n9528), .C1(
        pipeline_csr_mscratch[8]), .C2(n11268), .A(n10621), .ZN(n10631) );
  OAI22_X2 U11162 ( .A1(n13099), .A2(n6840), .B1(n9460), .B2(n10622), .ZN(
        n10623) );
  INV_X4 U11163 ( .A(ext_interrupts[0]), .ZN(n10625) );
  NAND4_X2 U11164 ( .A1(pipeline_inst_DX[29]), .A2(pipeline_inst_DX[28]), .A3(
        pipeline_imm_31_), .A4(pipeline_inst_DX[30]), .ZN(n13101) );
  INV_X4 U11165 ( .A(n13101), .ZN(n11111) );
  AOI221_X2 U11166 ( .B1(n6697), .B2(pipeline_csr_mie[8]), .C1(n11229), .C2(
        n10635), .A(n6818), .ZN(n10624) );
  OAI221_X2 U11167 ( .B1(n10625), .B2(n13103), .C1(n11997), .C2(n11262), .A(
        n10624), .ZN(n10628) );
  OAI22_X2 U11169 ( .A1(n1263), .A2(n11261), .B1(n1491), .B2(n13114), .ZN(
        n10626) );
  NOR3_X2 U11170 ( .A1(n10628), .A2(n10627), .A3(n10626), .ZN(n10629) );
  NOR2_X2 U11171 ( .A1(n6793), .A2(n10632), .ZN(n10633) );
  INV_X4 U11172 ( .A(n11999), .ZN(n12007) );
  NAND2_X2 U11173 ( .A1(n12007), .A2(n13130), .ZN(n10634) );
  MUX2_X2 U11174 ( .A(n10635), .B(n10634), .S(n6708), .Z(n6200) );
  OAI22_X2 U11175 ( .A1(n12007), .A2(n9516), .B1(n1523), .B2(n6660), .ZN(n6215) );
  INV_X4 U11176 ( .A(pipeline_md_N275), .ZN(n10636) );
  OAI22_X2 U11177 ( .A1(n1111), .A2(n9504), .B1(n12765), .B2(n10636), .ZN(
        n10637) );
  AOI221_X2 U11178 ( .B1(pipeline_md_N53), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[24]), .A(n10637), .ZN(n10638) );
  INV_X4 U11179 ( .A(n10638), .ZN(n5676) );
  INV_X4 U11180 ( .A(pipeline_md_result_muxed[56]), .ZN(n10640) );
  NOR2_X2 U11181 ( .A1(pipeline_md_N339), .A2(pipeline_md_resp_result[24]), 
        .ZN(n10639) );
  OAI22_X2 U11182 ( .A1(n10640), .A2(n6692), .B1(n10639), .B2(n6667), .ZN(
        n10641) );
  AOI221_X2 U11183 ( .B1(pipeline_md_N152), .B2(n6755), .C1(pipeline_md_N120), 
        .C2(n6754), .A(n10641), .ZN(n10644) );
  NOR2_X2 U11184 ( .A1(n1111), .A2(n6693), .ZN(n10642) );
  AOI221_X2 U11185 ( .B1(pipeline_md_N210), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[24]), .A(n10642), .ZN(n10643) );
  NAND2_X2 U11186 ( .A1(n10644), .A2(n10643), .ZN(n5629) );
  NAND2_X2 U11187 ( .A1(n11229), .A2(n10645), .ZN(n10646) );
  OAI221_X2 U11188 ( .B1(n1539), .B2(n9462), .C1(n11970), .C2(n9464), .A(
        n10646), .ZN(n10647) );
  AOI221_X2 U11189 ( .B1(n11138), .B2(n10648), .C1(n11136), .C2(
        ext_interrupts[16]), .A(n10647), .ZN(n10659) );
  OAI22_X2 U11190 ( .A1(n13111), .A2(n6876), .B1(n11269), .B2(n10649), .ZN(
        n10650) );
  AOI221_X2 U11191 ( .B1(n9527), .B2(n10651), .C1(pipeline_csr_mtime_full[24]), 
        .C2(n13108), .A(n10650), .ZN(n10658) );
  OAI22_X2 U11192 ( .A1(n13105), .A2(n6877), .B1(n11235), .B2(n10652), .ZN(
        n10653) );
  AOI221_X2 U11193 ( .B1(pipeline_csr_mscratch[24]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[24]), .C2(n13116), .A(n10653), .ZN(n10657) );
  OAI22_X2 U11194 ( .A1(n9460), .A2(n10654), .B1(n9526), .B2(n6833), .ZN(
        n10655) );
  AOI221_X2 U11195 ( .B1(pipeline_csr_cycle_full[56]), .B2(n11233), .C1(
        pipeline_csr_instret_full[56]), .C2(n11105), .A(n10655), .ZN(n10656)
         );
  NOR2_X2 U11196 ( .A1(pipeline_rs1_data_bypassed[24]), .A2(n9463), .ZN(n10660) );
  NOR2_X2 U11197 ( .A1(n6793), .A2(n10660), .ZN(n10662) );
  NAND2_X2 U11198 ( .A1(htif_pcr_req_data[24]), .A2(n13131), .ZN(n10661) );
  OAI221_X2 U11199 ( .B1(n7206), .B2(n10662), .C1(n12442), .C2(n9467), .A(
        n10661), .ZN(n11972) );
  INV_X4 U11200 ( .A(n11972), .ZN(n11982) );
  OAI22_X2 U11201 ( .A1(n11982), .A2(n6690), .B1(n1215), .B2(n6708), .ZN(n6184) );
  OAI22_X2 U11202 ( .A1(n11982), .A2(n9516), .B1(n1539), .B2(n6660), .ZN(n6231) );
  INV_X4 U11203 ( .A(imem_haddr[4]), .ZN(n10663) );
  OAI22_X2 U11204 ( .A1(n12525), .A2(n12632), .B1(n9493), .B2(n10663), .ZN(
        n5967) );
  OAI22_X2 U11205 ( .A1(n12525), .A2(n9496), .B1(n719), .B2(n6662), .ZN(n5931)
         );
  INV_X4 U11206 ( .A(pipeline_md_N258), .ZN(n10664) );
  OAI22_X2 U11207 ( .A1(n13048), .A2(n9504), .B1(n12765), .B2(n10664), .ZN(
        n10665) );
  INV_X4 U11208 ( .A(n10666), .ZN(n5659) );
  INV_X4 U11209 ( .A(pipeline_md_result_muxed[39]), .ZN(n10668) );
  NOR2_X2 U11210 ( .A1(pipeline_md_N322), .A2(pipeline_md_resp_result[7]), 
        .ZN(n10667) );
  OAI22_X2 U11211 ( .A1(n10668), .A2(n6692), .B1(n10667), .B2(n6667), .ZN(
        n10669) );
  AOI221_X2 U11212 ( .B1(pipeline_md_N135), .B2(n6755), .C1(pipeline_md_N103), 
        .C2(n6754), .A(n10669), .ZN(n10672) );
  NOR2_X2 U11213 ( .A1(n13048), .A2(n6693), .ZN(n10670) );
  AOI221_X2 U11214 ( .B1(pipeline_md_N193), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[7]), .A(n10670), .ZN(n10671) );
  NAND2_X2 U11215 ( .A1(n10672), .A2(n10671), .ZN(n5646) );
  NAND2_X2 U11216 ( .A1(n11229), .A2(n10673), .ZN(n10674) );
  OAI221_X2 U11217 ( .B1(n1522), .B2(n9462), .C1(n11890), .C2(n9464), .A(
        n10674), .ZN(n10675) );
  AOI221_X2 U11218 ( .B1(n11138), .B2(n10676), .C1(n11136), .C2(
        pipeline_csr_mip_7_), .A(n10675), .ZN(n10687) );
  OAI22_X2 U11219 ( .A1(n13111), .A2(n6841), .B1(n11269), .B2(n10677), .ZN(
        n10678) );
  AOI221_X2 U11220 ( .B1(n9527), .B2(n10679), .C1(pipeline_csr_mtime_full[7]), 
        .C2(n13108), .A(n10678), .ZN(n10686) );
  AOI221_X2 U11222 ( .B1(pipeline_csr_mscratch[7]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[7]), .C2(n13116), .A(n10681), .ZN(n10685) );
  OAI22_X2 U11223 ( .A1(n9460), .A2(n10682), .B1(n9526), .B2(n6842), .ZN(
        n10683) );
  AOI221_X2 U11224 ( .B1(pipeline_csr_time_full[39]), .B2(n11257), .C1(
        pipeline_csr_instret_full[39]), .C2(n11105), .A(n10683), .ZN(n10684)
         );
  NOR2_X2 U11225 ( .A1(n6793), .A2(n10688), .ZN(n10689) );
  OAI22_X2 U11226 ( .A1(n11943), .A2(n6690), .B1(n1198), .B2(n6708), .ZN(n6201) );
  OAI22_X2 U11227 ( .A1(n11943), .A2(n9516), .B1(n1522), .B2(n6660), .ZN(n6214) );
  INV_X4 U11228 ( .A(pipeline_md_N274), .ZN(n10690) );
  OAI22_X2 U11229 ( .A1(n13066), .A2(n9504), .B1(n12765), .B2(n10690), .ZN(
        n10691) );
  AOI221_X2 U11230 ( .B1(pipeline_md_N52), .B2(n6798), .C1(n6808), .C2(n6979), 
        .A(n10691), .ZN(n10692) );
  INV_X4 U11231 ( .A(n10692), .ZN(n5675) );
  INV_X4 U11232 ( .A(pipeline_md_result_muxed[55]), .ZN(n10694) );
  NOR2_X2 U11233 ( .A1(pipeline_md_N338), .A2(pipeline_md_resp_result[23]), 
        .ZN(n10693) );
  OAI22_X2 U11234 ( .A1(n10694), .A2(n6692), .B1(n10693), .B2(n6667), .ZN(
        n10695) );
  AOI221_X2 U11235 ( .B1(pipeline_md_N151), .B2(n6755), .C1(pipeline_md_N119), 
        .C2(n6754), .A(n10695), .ZN(n10698) );
  NOR2_X2 U11236 ( .A1(n13066), .A2(n6693), .ZN(n10696) );
  AOI221_X2 U11237 ( .B1(pipeline_md_N209), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[23]), .A(n10696), .ZN(n10697) );
  NAND2_X2 U11238 ( .A1(n10698), .A2(n10697), .ZN(n5630) );
  NAND2_X2 U11239 ( .A1(n11229), .A2(n10699), .ZN(n10700) );
  OAI221_X2 U11240 ( .B1(n1538), .B2(n9462), .C1(n11855), .C2(n9464), .A(
        n10700), .ZN(n10701) );
  AOI221_X2 U11241 ( .B1(n11138), .B2(n10702), .C1(n11136), .C2(
        ext_interrupts[15]), .A(n10701), .ZN(n10713) );
  OAI22_X2 U11242 ( .A1(n13111), .A2(n6878), .B1(n11269), .B2(n10703), .ZN(
        n10704) );
  AOI221_X2 U11243 ( .B1(n9527), .B2(n10705), .C1(pipeline_csr_mtime_full[23]), 
        .C2(n13108), .A(n10704), .ZN(n10712) );
  OAI22_X2 U11244 ( .A1(n13105), .A2(n6879), .B1(n11235), .B2(n10706), .ZN(
        n10707) );
  AOI221_X2 U11245 ( .B1(pipeline_csr_mscratch[23]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[23]), .C2(n13116), .A(n10707), .ZN(n10711) );
  OAI22_X2 U11246 ( .A1(n9460), .A2(n10708), .B1(n9526), .B2(n6900), .ZN(
        n10709) );
  AOI221_X2 U11247 ( .B1(pipeline_csr_cycle_full[55]), .B2(n11233), .C1(
        pipeline_csr_instret_full[55]), .C2(n11105), .A(n10709), .ZN(n10710)
         );
  NOR2_X2 U11248 ( .A1(n6979), .A2(n9463), .ZN(n10714) );
  NOR2_X2 U11249 ( .A1(n6793), .A2(n10714), .ZN(n10716) );
  NAND2_X2 U11250 ( .A1(htif_pcr_req_data[23]), .A2(n13131), .ZN(n10715) );
  OAI221_X2 U11251 ( .B1(n7205), .B2(n10716), .C1(n12446), .C2(n9467), .A(
        n10715), .ZN(n11857) );
  INV_X4 U11252 ( .A(n11857), .ZN(n11867) );
  OAI22_X2 U11253 ( .A1(n11867), .A2(n6690), .B1(n1214), .B2(n6708), .ZN(n6185) );
  OAI22_X2 U11254 ( .A1(n11867), .A2(n9516), .B1(n1538), .B2(n6660), .ZN(n6230) );
  INV_X4 U11255 ( .A(pipeline_md_N257), .ZN(n10717) );
  OAI22_X2 U11256 ( .A1(n13049), .A2(n9504), .B1(n12765), .B2(n10717), .ZN(
        n10718) );
  INV_X4 U11257 ( .A(n10719), .ZN(n5658) );
  INV_X4 U11258 ( .A(pipeline_md_result_muxed[38]), .ZN(n10721) );
  NOR2_X2 U11259 ( .A1(pipeline_md_N321), .A2(pipeline_md_resp_result[6]), 
        .ZN(n10720) );
  OAI22_X2 U11260 ( .A1(n10721), .A2(n6692), .B1(n10720), .B2(n6667), .ZN(
        n10722) );
  AOI221_X2 U11261 ( .B1(pipeline_md_N134), .B2(n6755), .C1(pipeline_md_N102), 
        .C2(n6754), .A(n10722), .ZN(n10725) );
  NOR2_X2 U11262 ( .A1(n13049), .A2(n6693), .ZN(n10723) );
  AOI221_X2 U11263 ( .B1(pipeline_md_N192), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[6]), .A(n10723), .ZN(n10724) );
  NAND2_X2 U11264 ( .A1(n10725), .A2(n10724), .ZN(n5647) );
  OAI22_X2 U11265 ( .A1(n1489), .A2(n13114), .B1(n11814), .B2(n11262), .ZN(
        n10726) );
  AOI221_X2 U11266 ( .B1(n11229), .B2(pipeline_csr_mtvec[6]), .C1(n6697), .C2(
        n10727), .A(n10726), .ZN(n10738) );
  OAI22_X2 U11267 ( .A1(n1389), .A2(n9460), .B1(n1160), .B2(n13099), .ZN(
        n10728) );
  AOI221_X2 U11268 ( .B1(n9527), .B2(n10730), .C1(n9461), .C2(n10729), .A(
        n10728), .ZN(n10737) );
  OAI22_X2 U11269 ( .A1(n11269), .A2(n10731), .B1(n11264), .B2(n6824), .ZN(
        n10732) );
  AOI221_X2 U11270 ( .B1(pipeline_csr_mtime_full[38]), .B2(n9528), .C1(
        pipeline_csr_mscratch[6]), .C2(n11268), .A(n10732), .ZN(n10736) );
  OAI22_X2 U11271 ( .A1(n13105), .A2(n6913), .B1(n13098), .B2(n10733), .ZN(
        n10734) );
  NOR2_X2 U11272 ( .A1(n6793), .A2(n10739), .ZN(n10740) );
  OAI221_X2 U11273 ( .B1(n7186), .B2(n10740), .C1(n12513), .C2(n9467), .A(
        n3715), .ZN(n11816) );
  INV_X4 U11274 ( .A(n11816), .ZN(n11824) );
  OAI22_X2 U11275 ( .A1(n11824), .A2(n6690), .B1(n1197), .B2(n6708), .ZN(n6202) );
  OAI22_X2 U11276 ( .A1(n11824), .A2(n9516), .B1(n1521), .B2(n6660), .ZN(n6213) );
  INV_X4 U11277 ( .A(pipeline_md_N273), .ZN(n10741) );
  OAI22_X2 U11278 ( .A1(n13067), .A2(n9504), .B1(n9505), .B2(n10741), .ZN(
        n10742) );
  AOI221_X2 U11279 ( .B1(pipeline_md_N51), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[22]), .A(n10742), .ZN(n10743) );
  INV_X4 U11280 ( .A(n10743), .ZN(n5674) );
  INV_X4 U11281 ( .A(pipeline_md_result_muxed[54]), .ZN(n10745) );
  NOR2_X2 U11282 ( .A1(pipeline_md_N337), .A2(pipeline_md_resp_result[22]), 
        .ZN(n10744) );
  OAI22_X2 U11283 ( .A1(n10745), .A2(n6692), .B1(n10744), .B2(n6667), .ZN(
        n10746) );
  AOI221_X2 U11284 ( .B1(pipeline_md_N150), .B2(n6755), .C1(pipeline_md_N118), 
        .C2(n6754), .A(n10746), .ZN(n10749) );
  NOR2_X2 U11285 ( .A1(n13067), .A2(n6693), .ZN(n10747) );
  AOI221_X2 U11286 ( .B1(pipeline_md_N208), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[22]), .A(n10747), .ZN(n10748) );
  NAND2_X2 U11287 ( .A1(n10749), .A2(n10748), .ZN(n5631) );
  NAND2_X2 U11288 ( .A1(n11229), .A2(n10750), .ZN(n10751) );
  OAI221_X2 U11289 ( .B1(n1537), .B2(n9462), .C1(n11785), .C2(n9464), .A(
        n10751), .ZN(n10752) );
  AOI221_X2 U11290 ( .B1(n11138), .B2(n10753), .C1(n11136), .C2(
        ext_interrupts[14]), .A(n10752), .ZN(n10765) );
  AOI221_X2 U11291 ( .B1(n9527), .B2(n10756), .C1(pipeline_csr_mtime_full[22]), 
        .C2(n13108), .A(n10755), .ZN(n10764) );
  OAI22_X2 U11292 ( .A1(n13098), .A2(n10758), .B1(n11235), .B2(n10757), .ZN(
        n10759) );
  AOI221_X2 U11293 ( .B1(pipeline_csr_mscratch[22]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[22]), .C2(n13116), .A(n10759), .ZN(n10763) );
  OAI22_X2 U11294 ( .A1(n9526), .A2(n6863), .B1(n9460), .B2(n10760), .ZN(
        n10761) );
  AOI221_X2 U11295 ( .B1(pipeline_csr_time_full[54]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[54]), .C2(n11233), .A(n10761), .ZN(n10762) );
  NOR2_X2 U11296 ( .A1(pipeline_rs1_data_bypassed[22]), .A2(n9463), .ZN(n10766) );
  NOR2_X2 U11297 ( .A1(n6793), .A2(n10766), .ZN(n10767) );
  OAI221_X2 U11298 ( .B1(n7204), .B2(n10767), .C1(n12450), .C2(n9467), .A(
        n3760), .ZN(n11787) );
  INV_X4 U11299 ( .A(n11787), .ZN(n11795) );
  OAI22_X2 U11300 ( .A1(n11795), .A2(n6690), .B1(n1213), .B2(n6708), .ZN(n6186) );
  OAI22_X2 U11301 ( .A1(n11795), .A2(n9516), .B1(n1537), .B2(n6660), .ZN(n6229) );
  INV_X4 U11302 ( .A(pipeline_md_N256), .ZN(n10768) );
  OAI22_X2 U11303 ( .A1(n1092), .A2(n9504), .B1(n9505), .B2(n10768), .ZN(
        n10769) );
  INV_X4 U11304 ( .A(n10770), .ZN(n5657) );
  INV_X4 U11305 ( .A(pipeline_md_result_muxed[37]), .ZN(n10772) );
  NOR2_X2 U11306 ( .A1(pipeline_md_N320), .A2(pipeline_md_resp_result[5]), 
        .ZN(n10771) );
  OAI22_X2 U11307 ( .A1(n10772), .A2(n6692), .B1(n10771), .B2(n6667), .ZN(
        n10773) );
  AOI221_X2 U11308 ( .B1(pipeline_md_N133), .B2(n6755), .C1(pipeline_md_N101), 
        .C2(n6754), .A(n10773), .ZN(n10776) );
  NOR2_X2 U11309 ( .A1(n1092), .A2(n6693), .ZN(n10774) );
  AOI221_X2 U11310 ( .B1(pipeline_md_N191), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[5]), .A(n10774), .ZN(n10775) );
  NAND2_X2 U11311 ( .A1(n10776), .A2(n10775), .ZN(n5648) );
  NAND3_X2 U11312 ( .A1(n6843), .A2(n7075), .A3(n6664), .ZN(n10777) );
  NAND2_X2 U11313 ( .A1(n9466), .A2(pipeline_csr_mtimecmp[5]), .ZN(n10778) );
  OAI221_X2 U11314 ( .B1(n1520), .B2(n9462), .C1(n1166), .C2(n13113), .A(
        n10778), .ZN(n10779) );
  AOI221_X2 U11315 ( .B1(n11138), .B2(n10781), .C1(n9527), .C2(n10780), .A(
        n10779), .ZN(n10790) );
  OAI22_X2 U11316 ( .A1(n13112), .A2(n12821), .B1(n11737), .B2(n11262), .ZN(
        n10782) );
  OAI22_X2 U11317 ( .A1(n10783), .A2(n6890), .B1(n11264), .B2(n6751), .ZN(
        n10784) );
  AOI221_X2 U11318 ( .B1(pipeline_csr_from_host[5]), .B2(n9461), .C1(
        pipeline_csr_instret_full[37]), .C2(n11105), .A(n10784), .ZN(n10788)
         );
  OAI22_X2 U11319 ( .A1(n9526), .A2(n6891), .B1(n9460), .B2(n10785), .ZN(
        n10786) );
  AOI221_X2 U11320 ( .B1(pipeline_csr_time_full[37]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[37]), .C2(n11233), .A(n10786), .ZN(n10787) );
  NOR2_X2 U11321 ( .A1(n6793), .A2(n10791), .ZN(n10792) );
  OAI221_X2 U11322 ( .B1(n6816), .B2(n10792), .C1(n12517), .C2(n9467), .A(
        n3711), .ZN(n11739) );
  OAI22_X2 U11323 ( .A1(n6702), .A2(n11752), .B1(n1292), .B2(n9529), .ZN(n6171) );
  OAI22_X2 U11324 ( .A1(n11752), .A2(n9516), .B1(n1520), .B2(n6660), .ZN(n6212) );
  NAND2_X2 U11325 ( .A1(n10793), .A2(n13130), .ZN(n3689) );
  OAI22_X2 U11326 ( .A1(n6688), .A2(n11752), .B1(n1166), .B2(n9530), .ZN(n6139) );
  MUX2_X2 U11327 ( .A(n12597), .B(pipeline_PC_DX[31]), .S(n9522), .Z(n5876) );
  MUX2_X2 U11328 ( .A(n10794), .B(pipeline_PC_DX[30]), .S(n9524), .Z(n5878) );
  MUX2_X2 U11329 ( .A(n10795), .B(pipeline_PC_DX[29]), .S(n9522), .Z(n5880) );
  MUX2_X2 U11330 ( .A(n10796), .B(pipeline_PC_DX[28]), .S(n9524), .Z(n5882) );
  OAI22_X2 U11331 ( .A1(n12433), .A2(n12632), .B1(n9493), .B2(n9378), .ZN(
        n5944) );
  OAI22_X2 U11332 ( .A1(n12433), .A2(n9496), .B1(n742), .B2(n6662), .ZN(n5885)
         );
  MUX2_X2 U11333 ( .A(n10797), .B(pipeline_PC_DX[27]), .S(n9522), .Z(n5884) );
  INV_X4 U11334 ( .A(n13165), .ZN(n10798) );
  OAI22_X2 U11335 ( .A1(n12437), .A2(n9494), .B1(n9493), .B2(n10798), .ZN(
        n5945) );
  OAI22_X2 U11336 ( .A1(n12437), .A2(n9496), .B1(n741), .B2(n6662), .ZN(n5887)
         );
  MUX2_X2 U11337 ( .A(n10799), .B(pipeline_PC_DX[26]), .S(n9523), .Z(n5886) );
  OAI22_X2 U11338 ( .A1(n12441), .A2(n9494), .B1(n9493), .B2(n9364), .ZN(n5946) );
  OAI22_X2 U11339 ( .A1(n12441), .A2(n9496), .B1(n740), .B2(n6662), .ZN(n5889)
         );
  MUX2_X2 U11340 ( .A(n10800), .B(pipeline_PC_DX[25]), .S(n9522), .Z(n5888) );
  OAI22_X2 U11341 ( .A1(n12445), .A2(n12632), .B1(n9370), .B2(n9493), .ZN(
        n5947) );
  OAI22_X2 U11342 ( .A1(n12445), .A2(n9496), .B1(n739), .B2(n6662), .ZN(n5891)
         );
  MUX2_X2 U11343 ( .A(n10801), .B(pipeline_PC_DX[24]), .S(n9523), .Z(n5890) );
  OAI22_X2 U11344 ( .A1(n12449), .A2(n9496), .B1(n738), .B2(n6662), .ZN(n5893)
         );
  MUX2_X2 U11345 ( .A(n10802), .B(pipeline_PC_DX[23]), .S(n9522), .Z(n5892) );
  OAI22_X2 U11346 ( .A1(n12453), .A2(n9494), .B1(n9493), .B2(n9366), .ZN(n5949) );
  OAI22_X2 U11347 ( .A1(n12453), .A2(n9496), .B1(n737), .B2(n6662), .ZN(n5895)
         );
  MUX2_X2 U11348 ( .A(n10803), .B(pipeline_PC_DX[22]), .S(n9525), .Z(n5894) );
  OAI22_X2 U11349 ( .A1(n12457), .A2(n12632), .B1(n9493), .B2(n9376), .ZN(
        n5950) );
  OAI22_X2 U11350 ( .A1(n12457), .A2(n9496), .B1(n736), .B2(n6662), .ZN(n5897)
         );
  MUX2_X2 U11351 ( .A(n10804), .B(pipeline_PC_DX[21]), .S(n9524), .Z(n5896) );
  OAI22_X2 U11352 ( .A1(n12461), .A2(n12632), .B1(n9493), .B2(n9368), .ZN(
        n5951) );
  OAI22_X2 U11353 ( .A1(n12461), .A2(n9497), .B1(n735), .B2(n6662), .ZN(n5899)
         );
  MUX2_X2 U11354 ( .A(n10805), .B(pipeline_PC_DX[20]), .S(n9523), .Z(n5898) );
  OAI22_X2 U11355 ( .A1(n12465), .A2(n12632), .B1(n9493), .B2(n9362), .ZN(
        n5952) );
  OAI22_X2 U11356 ( .A1(n12465), .A2(n9497), .B1(n734), .B2(n6662), .ZN(n5901)
         );
  MUX2_X2 U11357 ( .A(n10806), .B(pipeline_PC_DX[19]), .S(n9522), .Z(n5900) );
  OAI22_X2 U11358 ( .A1(n12469), .A2(n12632), .B1(n9493), .B2(n9374), .ZN(
        n5953) );
  OAI22_X2 U11359 ( .A1(n12469), .A2(n9497), .B1(n733), .B2(n6662), .ZN(n5903)
         );
  MUX2_X2 U11360 ( .A(n10807), .B(pipeline_PC_DX[18]), .S(n9524), .Z(n5902) );
  OAI22_X2 U11361 ( .A1(n12473), .A2(n12632), .B1(n9493), .B2(n10808), .ZN(
        n5954) );
  OAI22_X2 U11362 ( .A1(n12473), .A2(n9497), .B1(n732), .B2(n6662), .ZN(n5905)
         );
  MUX2_X2 U11363 ( .A(n10809), .B(pipeline_PC_DX[17]), .S(n9523), .Z(n5904) );
  OAI22_X2 U11364 ( .A1(n12476), .A2(n12632), .B1(n9493), .B2(n9346), .ZN(
        n5955) );
  OAI22_X2 U11365 ( .A1(n12476), .A2(n9497), .B1(n731), .B2(n6662), .ZN(n5907)
         );
  MUX2_X2 U11366 ( .A(n10810), .B(pipeline_PC_DX[16]), .S(n9525), .Z(n5906) );
  OAI22_X2 U11367 ( .A1(n12480), .A2(n12632), .B1(n9493), .B2(n9348), .ZN(
        n5956) );
  OAI22_X2 U11368 ( .A1(n12480), .A2(n9497), .B1(n730), .B2(n6662), .ZN(n5909)
         );
  MUX2_X2 U11369 ( .A(n10811), .B(pipeline_PC_DX[15]), .S(n9525), .Z(n5908) );
  OAI22_X2 U11370 ( .A1(n12484), .A2(n9494), .B1(n9493), .B2(n9350), .ZN(n5957) );
  OAI22_X2 U11371 ( .A1(n12484), .A2(n9497), .B1(n729), .B2(n6662), .ZN(n5911)
         );
  MUX2_X2 U11372 ( .A(n10812), .B(pipeline_PC_DX[14]), .S(n9524), .Z(n5910) );
  OAI22_X2 U11373 ( .A1(n12488), .A2(n9494), .B1(n9493), .B2(n9352), .ZN(n5958) );
  OAI22_X2 U11374 ( .A1(n12488), .A2(n9497), .B1(n728), .B2(n6662), .ZN(n5913)
         );
  MUX2_X2 U11375 ( .A(n10813), .B(pipeline_PC_DX[13]), .S(n9523), .Z(n5912) );
  OAI22_X2 U11376 ( .A1(n12492), .A2(n9497), .B1(n727), .B2(n6662), .ZN(n5915)
         );
  MUX2_X2 U11377 ( .A(n10814), .B(pipeline_PC_DX[12]), .S(n9522), .Z(n5914) );
  OAI22_X2 U11378 ( .A1(n12496), .A2(n9494), .B1(n9493), .B2(n9356), .ZN(n5960) );
  OAI22_X2 U11379 ( .A1(n12496), .A2(n9497), .B1(n726), .B2(n6662), .ZN(n5917)
         );
  MUX2_X2 U11380 ( .A(n10815), .B(pipeline_PC_DX[11]), .S(n9522), .Z(n5916) );
  OAI22_X2 U11381 ( .A1(n12500), .A2(n9497), .B1(n725), .B2(n6662), .ZN(n5919)
         );
  MUX2_X2 U11382 ( .A(n10816), .B(pipeline_PC_DX[10]), .S(n9524), .Z(n5918) );
  OAI221_X2 U11383 ( .B1(n12504), .B2(n9494), .C1(n9493), .C2(n9360), .A(
        n13130), .ZN(n5962) );
  OAI22_X2 U11384 ( .A1(n12504), .A2(n9497), .B1(n724), .B2(n6662), .ZN(n5921)
         );
  MUX2_X2 U11385 ( .A(n10817), .B(pipeline_PC_DX[9]), .S(n9522), .Z(n5920) );
  OAI22_X2 U11386 ( .A1(n12508), .A2(n9496), .B1(n723), .B2(n6662), .ZN(n5923)
         );
  MUX2_X2 U11387 ( .A(n10818), .B(pipeline_PC_DX[8]), .S(n9522), .Z(n5922) );
  OAI22_X2 U11388 ( .A1(n12512), .A2(n9494), .B1(n9493), .B2(n9344), .ZN(n5964) );
  OAI22_X2 U11389 ( .A1(n12512), .A2(n9497), .B1(n722), .B2(n6662), .ZN(n5925)
         );
  MUX2_X2 U11390 ( .A(n10819), .B(pipeline_PC_DX[7]), .S(n9522), .Z(n5924) );
  OAI22_X2 U11391 ( .A1(n12516), .A2(n9494), .B1(n9493), .B2(n9340), .ZN(n5965) );
  OAI22_X2 U11392 ( .A1(n12516), .A2(n9496), .B1(n721), .B2(n6662), .ZN(n5927)
         );
  MUX2_X2 U11393 ( .A(n10820), .B(pipeline_PC_DX[6]), .S(n9522), .Z(n5926) );
  INV_X4 U11394 ( .A(imem_haddr[5]), .ZN(n10821) );
  OAI22_X2 U11395 ( .A1(n12520), .A2(n9494), .B1(n9493), .B2(n10821), .ZN(
        n5966) );
  OAI22_X2 U11396 ( .A1(n12520), .A2(n9497), .B1(n720), .B2(n6662), .ZN(n5929)
         );
  MUX2_X2 U11397 ( .A(n10822), .B(pipeline_PC_DX[5]), .S(n9522), .Z(n5928) );
  MUX2_X2 U11398 ( .A(n12808), .B(pipeline_PC_DX[4]), .S(n9522), .Z(n5930) );
  MUX2_X2 U11399 ( .A(n12144), .B(pipeline_PC_DX[3]), .S(n9522), .Z(n5932) );
  MUX2_X2 U11400 ( .A(n12290), .B(pipeline_PC_DX[2]), .S(n9525), .Z(n5934) );
  NAND2_X2 U11401 ( .A1(pipeline_csr_N306), .A2(n6750), .ZN(n10823) );
  OAI221_X2 U11402 ( .B1(n11752), .B2(n6705), .C1(n1488), .C2(n6687), .A(
        n10823), .ZN(n5870) );
  OAI22_X2 U11403 ( .A1(n6659), .A2(n11752), .B1(n1260), .B2(n6689), .ZN(n6086) );
  INV_X4 U11404 ( .A(pipeline_md_N272), .ZN(n10826) );
  OAI22_X2 U11405 ( .A1(n1108), .A2(n9504), .B1(n12765), .B2(n10826), .ZN(
        n10827) );
  AOI221_X2 U11406 ( .B1(pipeline_md_N50), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[21]), .A(n10827), .ZN(n10828) );
  INV_X4 U11407 ( .A(n10828), .ZN(n5673) );
  INV_X4 U11408 ( .A(pipeline_md_result_muxed[53]), .ZN(n10830) );
  NOR2_X2 U11409 ( .A1(pipeline_md_N336), .A2(pipeline_md_resp_result[21]), 
        .ZN(n10829) );
  OAI22_X2 U11410 ( .A1(n10830), .A2(n6692), .B1(n10829), .B2(n6667), .ZN(
        n10831) );
  AOI221_X2 U11411 ( .B1(pipeline_md_N149), .B2(n6755), .C1(pipeline_md_N117), 
        .C2(n6754), .A(n10831), .ZN(n10834) );
  NOR2_X2 U11412 ( .A1(n1108), .A2(n6693), .ZN(n10832) );
  AOI221_X2 U11413 ( .B1(pipeline_md_N207), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[21]), .A(n10832), .ZN(n10833) );
  NAND2_X2 U11414 ( .A1(n10834), .A2(n10833), .ZN(n5632) );
  NAND2_X2 U11415 ( .A1(n11229), .A2(n10835), .ZN(n10836) );
  OAI221_X2 U11416 ( .B1(n1536), .B2(n9462), .C1(n11701), .C2(n9464), .A(
        n10836), .ZN(n10837) );
  AOI221_X2 U11417 ( .B1(n11138), .B2(n10838), .C1(n11136), .C2(
        ext_interrupts[13]), .A(n10837), .ZN(n10850) );
  AOI221_X2 U11418 ( .B1(n9527), .B2(n10841), .C1(pipeline_csr_mtime_full[21]), 
        .C2(n13108), .A(n10840), .ZN(n10849) );
  OAI22_X2 U11419 ( .A1(n13098), .A2(n10843), .B1(n11235), .B2(n10842), .ZN(
        n10844) );
  AOI221_X2 U11420 ( .B1(pipeline_csr_mscratch[21]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[21]), .C2(n13116), .A(n10844), .ZN(n10848) );
  OAI22_X2 U11421 ( .A1(n9526), .A2(n6892), .B1(n9460), .B2(n10845), .ZN(
        n10846) );
  AOI221_X2 U11422 ( .B1(pipeline_csr_time_full[53]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[53]), .C2(n11233), .A(n10846), .ZN(n10847) );
  NOR2_X2 U11423 ( .A1(pipeline_rs1_data_bypassed[21]), .A2(n9463), .ZN(n10851) );
  NOR2_X2 U11424 ( .A1(n6793), .A2(n10851), .ZN(n10852) );
  OAI221_X2 U11425 ( .B1(n7203), .B2(n10852), .C1(n12454), .C2(n9467), .A(
        n3757), .ZN(n11703) );
  INV_X4 U11426 ( .A(n11703), .ZN(n11711) );
  OAI22_X2 U11427 ( .A1(n11711), .A2(n6690), .B1(n1212), .B2(n6708), .ZN(n6187) );
  OAI22_X2 U11428 ( .A1(n11711), .A2(n9516), .B1(n1536), .B2(n6660), .ZN(n6228) );
  INV_X4 U11429 ( .A(pipeline_md_N263), .ZN(n10853) );
  OAI22_X2 U11430 ( .A1(n1099), .A2(n9504), .B1(n9505), .B2(n10853), .ZN(
        n10854) );
  INV_X4 U11431 ( .A(n10855), .ZN(n5664) );
  INV_X4 U11432 ( .A(pipeline_md_result_muxed[44]), .ZN(n10857) );
  NOR2_X2 U11433 ( .A1(pipeline_md_N327), .A2(pipeline_md_resp_result[12]), 
        .ZN(n10856) );
  OAI22_X2 U11434 ( .A1(n10857), .A2(n6692), .B1(n10856), .B2(n6667), .ZN(
        n10858) );
  AOI221_X2 U11435 ( .B1(pipeline_md_N140), .B2(n6755), .C1(pipeline_md_N108), 
        .C2(n6754), .A(n10858), .ZN(n10861) );
  NOR2_X2 U11436 ( .A1(n1099), .A2(n6693), .ZN(n10859) );
  AOI221_X2 U11437 ( .B1(pipeline_md_N198), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[12]), .A(n10859), .ZN(n10860) );
  NAND2_X2 U11438 ( .A1(n10861), .A2(n10860), .ZN(n5641) );
  NAND2_X2 U11439 ( .A1(n11229), .A2(n10862), .ZN(n10863) );
  OAI221_X2 U11440 ( .B1(n1527), .B2(n9462), .C1(n11660), .C2(n9464), .A(
        n10863), .ZN(n10864) );
  AOI221_X2 U11441 ( .B1(n11138), .B2(n10865), .C1(n11136), .C2(
        ext_interrupts[4]), .A(n10864), .ZN(n10877) );
  AOI221_X2 U11442 ( .B1(n9527), .B2(n10868), .C1(pipeline_csr_mtime_full[12]), 
        .C2(n13108), .A(n10867), .ZN(n10876) );
  OAI22_X2 U11443 ( .A1(n13098), .A2(n10870), .B1(n11235), .B2(n10869), .ZN(
        n10871) );
  AOI221_X2 U11444 ( .B1(pipeline_csr_mscratch[12]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[12]), .C2(n13116), .A(n10871), .ZN(n10875) );
  OAI22_X2 U11445 ( .A1(n9526), .A2(n6883), .B1(n9460), .B2(n10872), .ZN(
        n10873) );
  AOI221_X2 U11446 ( .B1(pipeline_csr_time_full[44]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[44]), .C2(n11233), .A(n10873), .ZN(n10874) );
  NOR2_X2 U11447 ( .A1(n6793), .A2(n10878), .ZN(n10879) );
  OAI221_X2 U11448 ( .B1(n7199), .B2(n10879), .C1(n12489), .C2(n9467), .A(
        n3730), .ZN(n11662) );
  INV_X4 U11449 ( .A(n11662), .ZN(n11670) );
  OAI22_X2 U11450 ( .A1(n11670), .A2(n6690), .B1(n1203), .B2(n6708), .ZN(n6196) );
  OAI22_X2 U11451 ( .A1(n11670), .A2(n9516), .B1(n1527), .B2(n6660), .ZN(n6219) );
  INV_X4 U11452 ( .A(pipeline_md_N271), .ZN(n10880) );
  OAI22_X2 U11453 ( .A1(n1107), .A2(n9504), .B1(n12765), .B2(n10880), .ZN(
        n10881) );
  AOI221_X2 U11454 ( .B1(pipeline_md_N49), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[20]), .A(n10881), .ZN(n10882) );
  INV_X4 U11455 ( .A(n10882), .ZN(n5672) );
  INV_X4 U11456 ( .A(pipeline_md_result_muxed[52]), .ZN(n10884) );
  NOR2_X2 U11457 ( .A1(pipeline_md_N335), .A2(pipeline_md_resp_result[20]), 
        .ZN(n10883) );
  OAI22_X2 U11458 ( .A1(n10884), .A2(n6692), .B1(n10883), .B2(n6667), .ZN(
        n10885) );
  AOI221_X2 U11459 ( .B1(pipeline_md_N148), .B2(n6755), .C1(pipeline_md_N116), 
        .C2(n6754), .A(n10885), .ZN(n10888) );
  NOR2_X2 U11460 ( .A1(n1107), .A2(n6693), .ZN(n10886) );
  AOI221_X2 U11461 ( .B1(pipeline_md_N206), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[20]), .A(n10886), .ZN(n10887) );
  NAND2_X2 U11462 ( .A1(n10888), .A2(n10887), .ZN(n5633) );
  NAND2_X2 U11463 ( .A1(n11105), .A2(n10889), .ZN(n10890) );
  OAI221_X2 U11464 ( .B1(n11264), .B2(n6822), .C1(n11269), .C2(n10891), .A(
        n10890), .ZN(n10892) );
  AOI221_X2 U11465 ( .B1(pipeline_csr_mtime_full[52]), .B2(n9528), .C1(
        pipeline_csr_mscratch[20]), .C2(n11268), .A(n10892), .ZN(n10904) );
  OAI22_X2 U11466 ( .A1(n13099), .A2(n6880), .B1(n9460), .B2(n10893), .ZN(
        n10894) );
  INV_X4 U11467 ( .A(ext_interrupts[12]), .ZN(n10898) );
  AOI221_X2 U11468 ( .B1(n6697), .B2(n10896), .C1(n11229), .C2(n10895), .A(
        n6818), .ZN(n10897) );
  OAI221_X2 U11469 ( .B1(n10898), .B2(n13103), .C1(n11627), .C2(n9464), .A(
        n10897), .ZN(n10901) );
  OAI22_X2 U11471 ( .A1(n1275), .A2(n11261), .B1(n1503), .B2(n13114), .ZN(
        n10899) );
  NOR3_X2 U11472 ( .A1(n10901), .A2(n10900), .A3(n10899), .ZN(n10902) );
  NOR2_X2 U11473 ( .A1(pipeline_rs1_data_bypassed[20]), .A2(n9463), .ZN(n10905) );
  NOR2_X2 U11474 ( .A1(n6793), .A2(n10905), .ZN(n10906) );
  OAI221_X2 U11475 ( .B1(n7187), .B2(n10906), .C1(n12458), .C2(n9467), .A(
        n3754), .ZN(n11629) );
  INV_X4 U11476 ( .A(n11629), .ZN(n11637) );
  OAI22_X2 U11477 ( .A1(n11637), .A2(n6690), .B1(n1211), .B2(n6708), .ZN(n6188) );
  OAI22_X2 U11478 ( .A1(n11637), .A2(n9516), .B1(n1535), .B2(n6660), .ZN(n6227) );
  INV_X4 U11479 ( .A(pipeline_md_N262), .ZN(n10907) );
  OAI22_X2 U11480 ( .A1(n13036), .A2(n9504), .B1(n12765), .B2(n10907), .ZN(
        n10908) );
  INV_X4 U11481 ( .A(n10909), .ZN(n5663) );
  INV_X4 U11482 ( .A(pipeline_md_result_muxed[43]), .ZN(n10911) );
  NOR2_X2 U11483 ( .A1(pipeline_md_N326), .A2(pipeline_md_resp_result[11]), 
        .ZN(n10910) );
  OAI22_X2 U11484 ( .A1(n10911), .A2(n6692), .B1(n10910), .B2(n6667), .ZN(
        n10912) );
  AOI221_X2 U11485 ( .B1(pipeline_md_N139), .B2(n6755), .C1(pipeline_md_N107), 
        .C2(n6754), .A(n10912), .ZN(n10915) );
  NOR2_X2 U11486 ( .A1(n13036), .A2(n6693), .ZN(n10913) );
  AOI221_X2 U11487 ( .B1(pipeline_md_N197), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[11]), .A(n10913), .ZN(n10914) );
  NAND2_X2 U11488 ( .A1(n10915), .A2(n10914), .ZN(n5642) );
  NAND2_X2 U11489 ( .A1(n11229), .A2(n10916), .ZN(n10917) );
  OAI221_X2 U11490 ( .B1(n1526), .B2(n9462), .C1(n11593), .C2(n9464), .A(
        n10917), .ZN(n10918) );
  AOI221_X2 U11491 ( .B1(n11138), .B2(n10919), .C1(n11136), .C2(
        ext_interrupts[3]), .A(n10918), .ZN(n10931) );
  AOI221_X2 U11492 ( .B1(n9527), .B2(n10922), .C1(pipeline_csr_mtime_full[11]), 
        .C2(n13108), .A(n10921), .ZN(n10930) );
  OAI22_X2 U11493 ( .A1(n13098), .A2(n10924), .B1(n11235), .B2(n10923), .ZN(
        n10925) );
  AOI221_X2 U11494 ( .B1(pipeline_csr_mscratch[11]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[11]), .C2(n13116), .A(n10925), .ZN(n10929) );
  OAI22_X2 U11495 ( .A1(n9526), .A2(n6893), .B1(n9460), .B2(n10926), .ZN(
        n10927) );
  AOI221_X2 U11496 ( .B1(pipeline_csr_time_full[43]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[43]), .C2(n11233), .A(n10927), .ZN(n10928) );
  NOR2_X2 U11497 ( .A1(n6793), .A2(n10932), .ZN(n10933) );
  OAI221_X2 U11498 ( .B1(n7200), .B2(n10933), .C1(n12493), .C2(n9467), .A(
        n3727), .ZN(n11595) );
  INV_X4 U11499 ( .A(n11595), .ZN(n11603) );
  OAI22_X2 U11500 ( .A1(n11603), .A2(n6690), .B1(n1202), .B2(n6708), .ZN(n6197) );
  OAI22_X2 U11501 ( .A1(n11603), .A2(n9516), .B1(n1526), .B2(n6660), .ZN(n6218) );
  INV_X4 U11502 ( .A(pipeline_md_N270), .ZN(n10934) );
  OAI22_X2 U11503 ( .A1(n13063), .A2(n9504), .B1(n12765), .B2(n10934), .ZN(
        n10935) );
  AOI221_X2 U11504 ( .B1(pipeline_md_N48), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[19]), .A(n10935), .ZN(n10936) );
  INV_X4 U11505 ( .A(n10936), .ZN(n5671) );
  INV_X4 U11506 ( .A(pipeline_md_result_muxed[51]), .ZN(n10938) );
  NOR2_X2 U11507 ( .A1(pipeline_md_N334), .A2(pipeline_md_resp_result[19]), 
        .ZN(n10937) );
  OAI22_X2 U11508 ( .A1(n10938), .A2(n6692), .B1(n10937), .B2(n6667), .ZN(
        n10939) );
  AOI221_X2 U11509 ( .B1(pipeline_md_N147), .B2(n6755), .C1(pipeline_md_N115), 
        .C2(n6754), .A(n10939), .ZN(n10942) );
  NOR2_X2 U11510 ( .A1(n13063), .A2(n6693), .ZN(n10940) );
  AOI221_X2 U11511 ( .B1(pipeline_md_N205), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[19]), .A(n10940), .ZN(n10941) );
  NAND2_X2 U11512 ( .A1(n10942), .A2(n10941), .ZN(n5634) );
  NAND2_X2 U11513 ( .A1(n11229), .A2(n10943), .ZN(n10944) );
  OAI221_X2 U11514 ( .B1(n1534), .B2(n9462), .C1(n11555), .C2(n9464), .A(
        n10944), .ZN(n10945) );
  AOI221_X2 U11515 ( .B1(n11138), .B2(n10946), .C1(n11136), .C2(
        ext_interrupts[11]), .A(n10945), .ZN(n10958) );
  AOI221_X2 U11516 ( .B1(n9527), .B2(n10949), .C1(pipeline_csr_mtime_full[19]), 
        .C2(n13108), .A(n10948), .ZN(n10957) );
  OAI22_X2 U11517 ( .A1(n13098), .A2(n10951), .B1(n11235), .B2(n10950), .ZN(
        n10952) );
  AOI221_X2 U11518 ( .B1(pipeline_csr_mscratch[19]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[19]), .C2(n13116), .A(n10952), .ZN(n10956) );
  OAI22_X2 U11519 ( .A1(n9526), .A2(n6894), .B1(n9460), .B2(n10953), .ZN(
        n10954) );
  AOI221_X2 U11520 ( .B1(pipeline_csr_time_full[51]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[51]), .C2(n11233), .A(n10954), .ZN(n10955) );
  NOR2_X2 U11521 ( .A1(n6793), .A2(n10959), .ZN(n10960) );
  OAI221_X2 U11522 ( .B1(n7194), .B2(n10960), .C1(n12462), .C2(n9467), .A(
        n3751), .ZN(n11557) );
  INV_X4 U11523 ( .A(n11557), .ZN(n11565) );
  OAI22_X2 U11524 ( .A1(n11565), .A2(n6690), .B1(n1210), .B2(n6708), .ZN(n6189) );
  OAI22_X2 U11525 ( .A1(n11565), .A2(n9516), .B1(n1534), .B2(n6660), .ZN(n6226) );
  INV_X4 U11526 ( .A(pipeline_md_N261), .ZN(n10961) );
  OAI22_X2 U11527 ( .A1(n13037), .A2(n9504), .B1(n12765), .B2(n10961), .ZN(
        n10962) );
  INV_X4 U11528 ( .A(n10963), .ZN(n5662) );
  INV_X4 U11529 ( .A(pipeline_md_result_muxed[42]), .ZN(n10965) );
  NOR2_X2 U11530 ( .A1(pipeline_md_N325), .A2(pipeline_md_resp_result[10]), 
        .ZN(n10964) );
  OAI22_X2 U11531 ( .A1(n10965), .A2(n6692), .B1(n10964), .B2(n6667), .ZN(
        n10966) );
  AOI221_X2 U11532 ( .B1(pipeline_md_N138), .B2(n6755), .C1(pipeline_md_N106), 
        .C2(n6754), .A(n10966), .ZN(n10969) );
  NOR2_X2 U11533 ( .A1(n13037), .A2(n6693), .ZN(n10967) );
  AOI221_X2 U11534 ( .B1(pipeline_md_N196), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[10]), .A(n10967), .ZN(n10968) );
  NAND2_X2 U11535 ( .A1(n10969), .A2(n10968), .ZN(n5643) );
  NAND2_X2 U11536 ( .A1(n11229), .A2(n10970), .ZN(n10971) );
  OAI221_X2 U11537 ( .B1(n1525), .B2(n9462), .C1(n11517), .C2(n9464), .A(
        n10971), .ZN(n10972) );
  AOI221_X2 U11538 ( .B1(n11138), .B2(n10973), .C1(n11136), .C2(
        ext_interrupts[2]), .A(n10972), .ZN(n10985) );
  AOI221_X2 U11539 ( .B1(n9527), .B2(n10976), .C1(pipeline_csr_mtime_full[10]), 
        .C2(n13108), .A(n10975), .ZN(n10984) );
  OAI22_X2 U11540 ( .A1(n13098), .A2(n10978), .B1(n11235), .B2(n10977), .ZN(
        n10979) );
  AOI221_X2 U11541 ( .B1(pipeline_csr_mscratch[10]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[10]), .C2(n13116), .A(n10979), .ZN(n10983) );
  OAI22_X2 U11542 ( .A1(n9526), .A2(n6884), .B1(n9460), .B2(n10980), .ZN(
        n10981) );
  AOI221_X2 U11543 ( .B1(pipeline_csr_time_full[42]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[42]), .C2(n11233), .A(n10981), .ZN(n10982) );
  NOR2_X2 U11544 ( .A1(n6793), .A2(n10986), .ZN(n10987) );
  OAI221_X2 U11545 ( .B1(n7201), .B2(n10987), .C1(n12497), .C2(n9467), .A(
        n3724), .ZN(n11519) );
  INV_X4 U11546 ( .A(n11519), .ZN(n11527) );
  OAI22_X2 U11547 ( .A1(n11527), .A2(n6690), .B1(n1201), .B2(n6708), .ZN(n6198) );
  OAI22_X2 U11548 ( .A1(n11527), .A2(n9516), .B1(n1525), .B2(n6660), .ZN(n6217) );
  INV_X4 U11549 ( .A(pipeline_md_N269), .ZN(n10988) );
  OAI22_X2 U11550 ( .A1(n13064), .A2(n9504), .B1(n12765), .B2(n10988), .ZN(
        n10989) );
  AOI221_X2 U11551 ( .B1(pipeline_md_N47), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[18]), .A(n10989), .ZN(n10990) );
  INV_X4 U11552 ( .A(n10990), .ZN(n5670) );
  INV_X4 U11553 ( .A(pipeline_md_result_muxed[50]), .ZN(n10992) );
  NOR2_X2 U11554 ( .A1(pipeline_md_N333), .A2(pipeline_md_resp_result[18]), 
        .ZN(n10991) );
  OAI22_X2 U11555 ( .A1(n10992), .A2(n6692), .B1(n10991), .B2(n6667), .ZN(
        n10993) );
  AOI221_X2 U11556 ( .B1(pipeline_md_N146), .B2(n6755), .C1(pipeline_md_N114), 
        .C2(n6754), .A(n10993), .ZN(n10996) );
  NOR2_X2 U11557 ( .A1(n13064), .A2(n6693), .ZN(n10994) );
  AOI221_X2 U11558 ( .B1(pipeline_md_N204), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[18]), .A(n10994), .ZN(n10995) );
  NAND2_X2 U11559 ( .A1(n10996), .A2(n10995), .ZN(n5635) );
  AOI221_X2 U11561 ( .B1(pipeline_csr_mscratch[18]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[18]), .C2(n13116), .A(n10999), .ZN(n11011) );
  OAI22_X2 U11562 ( .A1(n9526), .A2(n6864), .B1(n9460), .B2(n11000), .ZN(
        n11001) );
  AOI221_X2 U11563 ( .B1(pipeline_csr_time_full[50]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[50]), .C2(n11233), .A(n11001), .ZN(n11010) );
  NOR2_X2 U11564 ( .A1(n11481), .A2(n11262), .ZN(n11002) );
  AOI221_X2 U11565 ( .B1(n11229), .B2(n11003), .C1(n6697), .C2(
        pipeline_csr_mie[18]), .A(n11002), .ZN(n11004) );
  OAI221_X2 U11566 ( .B1(n1501), .B2(n13114), .C1(n13137), .C2(n13103), .A(
        n11004), .ZN(n11008) );
  OAI22_X2 U11567 ( .A1(n13111), .A2(n6881), .B1(n11269), .B2(n11005), .ZN(
        n11007) );
  OAI22_X2 U11568 ( .A1(n11264), .A2(n6851), .B1(n1273), .B2(n11261), .ZN(
        n11006) );
  NOR3_X2 U11569 ( .A1(n11008), .A2(n11007), .A3(n11006), .ZN(n11009) );
  NOR2_X2 U11570 ( .A1(pipeline_rs1_data_bypassed[18]), .A2(n9463), .ZN(n11012) );
  NOR2_X2 U11571 ( .A1(n6793), .A2(n11012), .ZN(n11013) );
  OAI221_X2 U11572 ( .B1(n7188), .B2(n11013), .C1(n12466), .C2(n9467), .A(
        n3748), .ZN(n11483) );
  INV_X4 U11573 ( .A(n11483), .ZN(n11491) );
  OAI22_X2 U11574 ( .A1(n11491), .A2(n6690), .B1(n1209), .B2(n6708), .ZN(n6190) );
  OAI22_X2 U11575 ( .A1(n11491), .A2(n9516), .B1(n1533), .B2(n6660), .ZN(n6225) );
  INV_X4 U11576 ( .A(pipeline_md_N264), .ZN(n11014) );
  OAI22_X2 U11577 ( .A1(n1100), .A2(n9504), .B1(n12765), .B2(n11014), .ZN(
        n11015) );
  AOI221_X2 U11578 ( .B1(pipeline_md_N42), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[13]), .A(n11015), .ZN(n11016) );
  INV_X4 U11579 ( .A(n11016), .ZN(n5665) );
  INV_X4 U11580 ( .A(pipeline_md_result_muxed[45]), .ZN(n11018) );
  NOR2_X2 U11581 ( .A1(pipeline_md_N328), .A2(pipeline_md_resp_result[13]), 
        .ZN(n11017) );
  OAI22_X2 U11582 ( .A1(n11018), .A2(n6692), .B1(n11017), .B2(n6667), .ZN(
        n11019) );
  AOI221_X2 U11583 ( .B1(pipeline_md_N141), .B2(n6755), .C1(pipeline_md_N109), 
        .C2(n6754), .A(n11019), .ZN(n11022) );
  NOR2_X2 U11584 ( .A1(n1100), .A2(n6693), .ZN(n11020) );
  AOI221_X2 U11585 ( .B1(pipeline_md_N199), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[13]), .A(n11020), .ZN(n11021) );
  NAND2_X2 U11586 ( .A1(n11022), .A2(n11021), .ZN(n5640) );
  NAND2_X2 U11587 ( .A1(n11229), .A2(n11023), .ZN(n11024) );
  OAI221_X2 U11588 ( .B1(n1528), .B2(n9462), .C1(n11451), .C2(n9464), .A(
        n11024), .ZN(n11025) );
  AOI221_X2 U11589 ( .B1(n11138), .B2(n11026), .C1(n11136), .C2(
        ext_interrupts[5]), .A(n11025), .ZN(n11038) );
  AOI221_X2 U11590 ( .B1(n9527), .B2(n11029), .C1(pipeline_csr_mtime_full[13]), 
        .C2(n13108), .A(n11028), .ZN(n11037) );
  OAI22_X2 U11591 ( .A1(n13098), .A2(n11031), .B1(n11235), .B2(n11030), .ZN(
        n11032) );
  AOI221_X2 U11592 ( .B1(pipeline_csr_mscratch[13]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[13]), .C2(n13116), .A(n11032), .ZN(n11036) );
  OAI22_X2 U11593 ( .A1(n9526), .A2(n6895), .B1(n9460), .B2(n11033), .ZN(
        n11034) );
  AOI221_X2 U11594 ( .B1(pipeline_csr_time_full[45]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[45]), .C2(n11233), .A(n11034), .ZN(n11035) );
  NOR2_X2 U11595 ( .A1(pipeline_rs1_data_bypassed[13]), .A2(n9463), .ZN(n11039) );
  NOR2_X2 U11596 ( .A1(n6793), .A2(n11039), .ZN(n11040) );
  OAI221_X2 U11597 ( .B1(n7198), .B2(n11040), .C1(n12485), .C2(n9467), .A(
        n3733), .ZN(n11453) );
  INV_X4 U11598 ( .A(n11453), .ZN(n11461) );
  OAI22_X2 U11599 ( .A1(n11461), .A2(n6690), .B1(n1204), .B2(n6708), .ZN(n6195) );
  OAI22_X2 U11600 ( .A1(n11461), .A2(n9516), .B1(n1528), .B2(n6660), .ZN(n6220) );
  INV_X4 U11601 ( .A(pipeline_md_N268), .ZN(n11041) );
  OAI22_X2 U11602 ( .A1(n1104), .A2(n9504), .B1(n12765), .B2(n11041), .ZN(
        n11042) );
  AOI221_X2 U11603 ( .B1(pipeline_md_N46), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[17]), .A(n11042), .ZN(n11043) );
  INV_X4 U11604 ( .A(n11043), .ZN(n5669) );
  INV_X4 U11605 ( .A(pipeline_md_result_muxed[49]), .ZN(n11045) );
  NOR2_X2 U11606 ( .A1(pipeline_md_N332), .A2(pipeline_md_resp_result[17]), 
        .ZN(n11044) );
  OAI22_X2 U11607 ( .A1(n11045), .A2(n6692), .B1(n11044), .B2(n6667), .ZN(
        n11046) );
  AOI221_X2 U11608 ( .B1(pipeline_md_N145), .B2(n6755), .C1(pipeline_md_N113), 
        .C2(n6754), .A(n11046), .ZN(n11049) );
  NOR2_X2 U11609 ( .A1(n1104), .A2(n6693), .ZN(n11047) );
  AOI221_X2 U11610 ( .B1(pipeline_md_N203), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[17]), .A(n11047), .ZN(n11048) );
  NAND2_X2 U11611 ( .A1(n11049), .A2(n11048), .ZN(n5636) );
  NAND2_X2 U11612 ( .A1(n11229), .A2(n11050), .ZN(n11051) );
  OAI221_X2 U11613 ( .B1(n1532), .B2(n9462), .C1(n11421), .C2(n9464), .A(
        n11051), .ZN(n11052) );
  AOI221_X2 U11614 ( .B1(n11138), .B2(n11053), .C1(n11136), .C2(
        ext_interrupts[9]), .A(n11052), .ZN(n11065) );
  AOI221_X2 U11615 ( .B1(n9527), .B2(n11056), .C1(pipeline_csr_mtime_full[17]), 
        .C2(n13108), .A(n11055), .ZN(n11064) );
  OAI22_X2 U11616 ( .A1(n13098), .A2(n11058), .B1(n11235), .B2(n11057), .ZN(
        n11059) );
  AOI221_X2 U11617 ( .B1(pipeline_csr_mscratch[17]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[17]), .C2(n13116), .A(n11059), .ZN(n11063) );
  OAI22_X2 U11618 ( .A1(n9526), .A2(n6896), .B1(n9460), .B2(n11060), .ZN(
        n11061) );
  AOI221_X2 U11619 ( .B1(pipeline_csr_time_full[49]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[49]), .C2(n11233), .A(n11061), .ZN(n11062) );
  NOR2_X2 U11620 ( .A1(pipeline_rs1_data_bypassed[17]), .A2(n9463), .ZN(n11066) );
  NOR2_X2 U11621 ( .A1(n6793), .A2(n11066), .ZN(n11067) );
  OAI221_X2 U11622 ( .B1(n7195), .B2(n11067), .C1(n12470), .C2(n9467), .A(
        n3745), .ZN(n11423) );
  INV_X4 U11623 ( .A(n11423), .ZN(n11431) );
  OAI22_X2 U11624 ( .A1(n11431), .A2(n6690), .B1(n1208), .B2(n6708), .ZN(n6191) );
  OAI22_X2 U11625 ( .A1(n11431), .A2(n9516), .B1(n1532), .B2(n6660), .ZN(n6224) );
  INV_X4 U11626 ( .A(pipeline_md_N267), .ZN(n11068) );
  OAI22_X2 U11627 ( .A1(n1103), .A2(n9504), .B1(n12765), .B2(n11068), .ZN(
        n11069) );
  INV_X4 U11628 ( .A(n11070), .ZN(n5668) );
  INV_X4 U11629 ( .A(pipeline_md_result_muxed[48]), .ZN(n11072) );
  NOR2_X2 U11630 ( .A1(pipeline_md_N331), .A2(pipeline_md_resp_result[16]), 
        .ZN(n11071) );
  OAI22_X2 U11631 ( .A1(n11072), .A2(n6692), .B1(n11071), .B2(n6667), .ZN(
        n11073) );
  AOI221_X2 U11632 ( .B1(pipeline_md_N144), .B2(n6755), .C1(pipeline_md_N112), 
        .C2(n6754), .A(n11073), .ZN(n11076) );
  NOR2_X2 U11633 ( .A1(n1103), .A2(n6693), .ZN(n11074) );
  AOI221_X2 U11634 ( .B1(pipeline_md_N202), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[16]), .A(n11074), .ZN(n11075) );
  NAND2_X2 U11635 ( .A1(n11076), .A2(n11075), .ZN(n5637) );
  NAND2_X2 U11636 ( .A1(n11229), .A2(n11077), .ZN(n11078) );
  OAI221_X2 U11637 ( .B1(n1531), .B2(n9462), .C1(n11382), .C2(n9464), .A(
        n11078), .ZN(n11079) );
  AOI221_X2 U11638 ( .B1(n11138), .B2(n11080), .C1(n11136), .C2(
        ext_interrupts[8]), .A(n11079), .ZN(n11092) );
  AOI221_X2 U11639 ( .B1(n9527), .B2(n11083), .C1(pipeline_csr_mtime_full[16]), 
        .C2(n13108), .A(n11082), .ZN(n11091) );
  OAI22_X2 U11640 ( .A1(n13098), .A2(n11085), .B1(n11235), .B2(n11084), .ZN(
        n11086) );
  AOI221_X2 U11641 ( .B1(pipeline_csr_mscratch[16]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[16]), .C2(n13116), .A(n11086), .ZN(n11090) );
  OAI22_X2 U11642 ( .A1(n9526), .A2(n6885), .B1(n9460), .B2(n11087), .ZN(
        n11088) );
  AOI221_X2 U11643 ( .B1(pipeline_csr_time_full[48]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[48]), .C2(n11233), .A(n11088), .ZN(n11089) );
  NOR2_X2 U11644 ( .A1(n6793), .A2(n11093), .ZN(n11094) );
  OAI221_X2 U11645 ( .B1(n7196), .B2(n11094), .C1(n12474), .C2(n9467), .A(
        n3742), .ZN(n11384) );
  INV_X4 U11646 ( .A(n11384), .ZN(n11392) );
  OAI22_X2 U11647 ( .A1(n11392), .A2(n6690), .B1(n1207), .B2(n6708), .ZN(n6192) );
  OAI22_X2 U11648 ( .A1(n11392), .A2(n9516), .B1(n1531), .B2(n6660), .ZN(n6223) );
  INV_X4 U11649 ( .A(pipeline_md_N266), .ZN(n11095) );
  OAI22_X2 U11650 ( .A1(n13039), .A2(n9504), .B1(n12765), .B2(n11095), .ZN(
        n11096) );
  INV_X4 U11651 ( .A(n11097), .ZN(n5667) );
  INV_X4 U11652 ( .A(pipeline_md_result_muxed[47]), .ZN(n11099) );
  NOR2_X2 U11653 ( .A1(pipeline_md_N330), .A2(pipeline_md_resp_result[15]), 
        .ZN(n11098) );
  OAI22_X2 U11654 ( .A1(n11099), .A2(n6692), .B1(n11098), .B2(n6667), .ZN(
        n11100) );
  AOI221_X2 U11655 ( .B1(pipeline_md_N143), .B2(n6755), .C1(pipeline_md_N111), 
        .C2(n6754), .A(n11100), .ZN(n11103) );
  NOR2_X2 U11656 ( .A1(n13039), .A2(n6693), .ZN(n11101) );
  AOI221_X2 U11657 ( .B1(pipeline_md_N201), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[15]), .A(n11101), .ZN(n11102) );
  NAND2_X2 U11658 ( .A1(n11103), .A2(n11102), .ZN(n5638) );
  NAND2_X2 U11659 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  OAI221_X2 U11660 ( .B1(n11264), .B2(n6865), .C1(n11269), .C2(n11107), .A(
        n11106), .ZN(n11108) );
  AOI221_X2 U11661 ( .B1(pipeline_csr_mtime_full[47]), .B2(n9528), .C1(
        pipeline_csr_mscratch[15]), .C2(n11268), .A(n11108), .ZN(n11121) );
  OAI22_X2 U11662 ( .A1(n13099), .A2(n6882), .B1(n9460), .B2(n11109), .ZN(
        n11110) );
  NAND2_X2 U11663 ( .A1(n7077), .A2(n11111), .ZN(n13110) );
  INV_X4 U11664 ( .A(n13110), .ZN(n11112) );
  AOI221_X2 U11665 ( .B1(n6697), .B2(n11114), .C1(n11229), .C2(n11113), .A(
        n11112), .ZN(n11115) );
  OAI221_X2 U11666 ( .B1(n6959), .B2(n13103), .C1(n11352), .C2(n9464), .A(
        n11115), .ZN(n11118) );
  OAI22_X2 U11668 ( .A1(n1270), .A2(n11261), .B1(n1498), .B2(n13114), .ZN(
        n11116) );
  NOR3_X2 U11669 ( .A1(n11118), .A2(n11117), .A3(n11116), .ZN(n11119) );
  NOR2_X2 U11670 ( .A1(n6793), .A2(n11122), .ZN(n11123) );
  OAI221_X2 U11671 ( .B1(n7189), .B2(n11123), .C1(n12477), .C2(n9467), .A(
        n3739), .ZN(n11354) );
  INV_X4 U11672 ( .A(n11354), .ZN(n11362) );
  OAI22_X2 U11673 ( .A1(n11362), .A2(n6690), .B1(n1206), .B2(n6708), .ZN(n6193) );
  OAI22_X2 U11674 ( .A1(n11362), .A2(n9516), .B1(n1530), .B2(n6660), .ZN(n6222) );
  INV_X4 U11675 ( .A(pipeline_md_N265), .ZN(n11124) );
  OAI22_X2 U11676 ( .A1(n13040), .A2(n9504), .B1(n9505), .B2(n11124), .ZN(
        n11125) );
  AOI221_X2 U11677 ( .B1(pipeline_md_N43), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[14]), .A(n11125), .ZN(n11126) );
  INV_X4 U11678 ( .A(n11126), .ZN(n5666) );
  INV_X4 U11679 ( .A(pipeline_md_result_muxed[46]), .ZN(n11128) );
  NOR2_X2 U11680 ( .A1(pipeline_md_N329), .A2(pipeline_md_resp_result[14]), 
        .ZN(n11127) );
  OAI22_X2 U11681 ( .A1(n11128), .A2(n6692), .B1(n11127), .B2(n6667), .ZN(
        n11129) );
  AOI221_X2 U11682 ( .B1(pipeline_md_N142), .B2(n6755), .C1(pipeline_md_N110), 
        .C2(n6754), .A(n11129), .ZN(n11132) );
  NOR2_X2 U11683 ( .A1(n13040), .A2(n6693), .ZN(n11130) );
  AOI221_X2 U11684 ( .B1(pipeline_md_N200), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[14]), .A(n11130), .ZN(n11131) );
  NAND2_X2 U11685 ( .A1(n11132), .A2(n11131), .ZN(n5639) );
  NAND2_X2 U11686 ( .A1(n11229), .A2(n11133), .ZN(n11134) );
  OAI221_X2 U11687 ( .B1(n1529), .B2(n9462), .C1(n11194), .C2(n9464), .A(
        n11134), .ZN(n11135) );
  AOI221_X2 U11688 ( .B1(n11138), .B2(n11137), .C1(n11136), .C2(
        ext_interrupts[6]), .A(n11135), .ZN(n11150) );
  AOI221_X2 U11689 ( .B1(n9527), .B2(n11141), .C1(pipeline_csr_mtime_full[14]), 
        .C2(n13108), .A(n11140), .ZN(n11149) );
  OAI22_X2 U11690 ( .A1(n13098), .A2(n11143), .B1(n11235), .B2(n11142), .ZN(
        n11144) );
  AOI221_X2 U11691 ( .B1(pipeline_csr_mscratch[14]), .B2(n11268), .C1(
        pipeline_csr_cycle_full[14]), .C2(n13116), .A(n11144), .ZN(n11148) );
  OAI22_X2 U11692 ( .A1(n9526), .A2(n6886), .B1(n9460), .B2(n11145), .ZN(
        n11146) );
  AOI221_X2 U11693 ( .B1(pipeline_csr_time_full[46]), .B2(n11257), .C1(
        pipeline_csr_cycle_full[46]), .C2(n11233), .A(n11146), .ZN(n11147) );
  NOR2_X2 U11694 ( .A1(pipeline_rs1_data_bypassed[14]), .A2(n9463), .ZN(n11151) );
  NOR2_X2 U11695 ( .A1(n6793), .A2(n11151), .ZN(n11152) );
  OAI221_X2 U11696 ( .B1(n7197), .B2(n11152), .C1(n12481), .C2(n9467), .A(
        n3736), .ZN(n11218) );
  INV_X4 U11697 ( .A(n11218), .ZN(n11328) );
  OAI22_X2 U11698 ( .A1(n11328), .A2(n6690), .B1(n1205), .B2(n6708), .ZN(n6194) );
  OAI22_X2 U11699 ( .A1(n11328), .A2(n9516), .B1(n1529), .B2(n6660), .ZN(n6221) );
  NAND2_X2 U11700 ( .A1(n9479), .A2(n11174), .ZN(n11153) );
  NAND2_X2 U11701 ( .A1(n11153), .A2(n9512), .ZN(n11164) );
  INV_X4 U11702 ( .A(n12791), .ZN(n12567) );
  NAND2_X2 U11703 ( .A1(n12567), .A2(pipeline_alu_src_b[4]), .ZN(n11579) );
  INV_X4 U11704 ( .A(n11579), .ZN(n12062) );
  NAND2_X2 U11705 ( .A1(n9509), .A2(n7005), .ZN(n11641) );
  MUX2_X2 U11706 ( .A(n7006), .B(n6997), .S(n9489), .Z(n11770) );
  NAND2_X2 U11707 ( .A1(n9510), .A2(n11770), .ZN(n11154) );
  NAND2_X2 U11708 ( .A1(n11641), .A2(n11154), .ZN(n12634) );
  NAND2_X2 U11709 ( .A1(n9471), .A2(n6980), .ZN(n11961) );
  NAND2_X2 U11710 ( .A1(n12276), .A2(pipeline_alu_src_a[24]), .ZN(n12098) );
  NAND2_X2 U11711 ( .A1(n11869), .A2(n6608), .ZN(n12210) );
  NAND2_X2 U11712 ( .A1(n9489), .A2(n6626), .ZN(n11775) );
  NAND4_X2 U11713 ( .A1(n11961), .A2(n12098), .A3(n12210), .A4(n11775), .ZN(
        n11500) );
  NAND2_X2 U11714 ( .A1(n12276), .A2(n6564), .ZN(n12654) );
  NAND2_X2 U11715 ( .A1(n11869), .A2(pipeline_alu_src_a[29]), .ZN(n11155) );
  NAND2_X2 U11716 ( .A1(n9489), .A2(n6560), .ZN(n12096) );
  NAND4_X2 U11717 ( .A1(n12212), .A2(n12654), .A3(n11155), .A4(n12096), .ZN(
        n11495) );
  INV_X4 U11718 ( .A(n12281), .ZN(n11498) );
  NAND2_X2 U11719 ( .A1(n9471), .A2(pipeline_alu_src_a[19]), .ZN(n11620) );
  NAND2_X2 U11720 ( .A1(n12276), .A2(pipeline_alu_src_a[20]), .ZN(n11777) );
  NAND2_X2 U11721 ( .A1(n9489), .A2(pipeline_alu_src_a[18]), .ZN(n11157) );
  NAND2_X2 U11722 ( .A1(n11869), .A2(pipeline_alu_src_a[21]), .ZN(n11959) );
  NAND4_X2 U11723 ( .A1(n11620), .A2(n11777), .A3(n11157), .A4(n11959), .ZN(
        n11801) );
  INV_X4 U11724 ( .A(n11801), .ZN(n11471) );
  OAI22_X2 U11725 ( .A1(n11498), .A2(n12776), .B1(n11471), .B2(n9507), .ZN(
        n11158) );
  AOI221_X2 U11726 ( .B1(n9511), .B2(n11500), .C1(n12780), .C2(n11495), .A(
        n11158), .ZN(n11162) );
  MUX2_X2 U11727 ( .A(n7005), .B(n6997), .S(n11404), .Z(n11160) );
  NAND2_X2 U11728 ( .A1(n11160), .A2(n11405), .ZN(n11501) );
  INV_X4 U11729 ( .A(n12794), .ZN(n12199) );
  NAND2_X2 U11730 ( .A1(n12199), .A2(n6600), .ZN(n12058) );
  INV_X4 U11731 ( .A(n12058), .ZN(n11161) );
  NAND2_X2 U11732 ( .A1(n11161), .A2(n9510), .ZN(n11645) );
  OAI22_X2 U11733 ( .A1(n11162), .A2(n12772), .B1(n11501), .B2(n11645), .ZN(
        n11163) );
  AOI221_X2 U11734 ( .B1(n11164), .B2(pipeline_alu_src_a[14]), .C1(n12062), 
        .C2(n12634), .A(n11163), .ZN(n11177) );
  INV_X4 U11735 ( .A(n11755), .ZN(n11466) );
  NOR2_X2 U11736 ( .A1(n11869), .A2(n11166), .ZN(n11167) );
  OAI22_X2 U11737 ( .A1(n11758), .A2(n9509), .B1(n11757), .B2(n9507), .ZN(
        n11170) );
  AOI221_X2 U11738 ( .B1(n9511), .B2(n11466), .C1(n12780), .C2(n11507), .A(
        n11170), .ZN(n11171) );
  INV_X4 U11739 ( .A(n11171), .ZN(n12650) );
  MUX2_X2 U11740 ( .A(n12793), .B(n9479), .S(n11570), .Z(n11172) );
  NOR2_X2 U11741 ( .A1(n9513), .A2(n11172), .ZN(n11173) );
  OAI22_X2 U11742 ( .A1(n12785), .A2(n12650), .B1(n11174), .B2(n11173), .ZN(
        n11175) );
  AOI221_X2 U11743 ( .B1(pipeline_alu_N73), .B2(n6813), .C1(pipeline_alu_N267), 
        .C2(n6812), .A(n11175), .ZN(n11176) );
  NAND2_X2 U11744 ( .A1(n11177), .A2(n11176), .ZN(dmem_haddr[14]) );
  MUX2_X2 U11745 ( .A(pipeline_alu_out_WB[14]), .B(dmem_haddr[14]), .S(n9522), 
        .Z(n5830) );
  NAND2_X2 U11746 ( .A1(n12832), .A2(n6922), .ZN(n11181) );
  NAND3_X2 U11747 ( .A1(imem_hresp), .A2(imem_hready), .A3(n11178), .ZN(
        n11180) );
  OAI22_X2 U11748 ( .A1(n11181), .A2(n11180), .B1(n799), .B2(n11179), .ZN(
        n6300) );
  INV_X4 U11749 ( .A(n11187), .ZN(n11182) );
  NAND2_X2 U11750 ( .A1(n6844), .A2(n11182), .ZN(n11185) );
  NAND2_X2 U11751 ( .A1(n12827), .A2(pipeline_ctrl_prev_ex_code_WB[3]), .ZN(
        n11183) );
  NAND2_X2 U11752 ( .A1(n11185), .A2(n11183), .ZN(n5978) );
  NAND3_X2 U11753 ( .A1(n7075), .A2(n7177), .A3(n6844), .ZN(n11184) );
  OAI221_X2 U11754 ( .B1(n10323), .B2(n11185), .C1(n780), .C2(n9523), .A(
        n11184), .ZN(n5977) );
  NOR2_X2 U11755 ( .A1(n9525), .A2(n11191), .ZN(n5979) );
  INV_X4 U11756 ( .A(n11185), .ZN(n11186) );
  NAND2_X2 U11757 ( .A1(n11186), .A2(pipeline_ctrl_N82), .ZN(n11190) );
  NAND2_X2 U11758 ( .A1(n799), .A2(n11187), .ZN(n11188) );
  MUX2_X2 U11759 ( .A(n781), .B(n11188), .S(n9524), .Z(n11189) );
  NAND2_X2 U11760 ( .A1(n11190), .A2(n11189), .ZN(n5976) );
  NAND2_X2 U11761 ( .A1(n6369), .A2(n12806), .ZN(n12805) );
  NAND2_X2 U11762 ( .A1(n11191), .A2(pipeline_ctrl_had_ex_WB), .ZN(n12292) );
  NAND3_X2 U11763 ( .A1(n9515), .A2(n12806), .A3(n11192), .ZN(n12617) );
  INV_X4 U11764 ( .A(n11192), .ZN(n11193) );
  OAI22_X2 U11765 ( .A1(n9515), .A2(n11194), .B1(n549), .B2(n9498), .ZN(n11195) );
  AOI221_X2 U11766 ( .B1(n12668), .B2(n11218), .C1(pipeline_alu_out_WB[14]), 
        .C2(n12809), .A(n11195), .ZN(n11196) );
  INV_X4 U11767 ( .A(n11196), .ZN(n5798) );
  NAND2_X2 U11768 ( .A1(pipeline_csr_N315), .A2(n6750), .ZN(n11197) );
  OAI221_X2 U11769 ( .B1(n11328), .B2(n6705), .C1(n1497), .C2(n6687), .A(
        n11197), .ZN(n5861) );
  OAI22_X2 U11770 ( .A1(n6659), .A2(n11328), .B1(n1269), .B2(n6689), .ZN(n6095) );
  NOR2_X2 U11771 ( .A1(n11283), .A2(n11318), .ZN(n11200) );
  INV_X4 U11772 ( .A(n11284), .ZN(n11199) );
  INV_X4 U11773 ( .A(pipeline_csr_N903), .ZN(n11201) );
  OAI22_X2 U11774 ( .A1(n6669), .A2(n11201), .B1(n12603), .B2(n11282), .ZN(
        pipeline_csr_N2164) );
  INV_X4 U11775 ( .A(pipeline_csr_N902), .ZN(n11202) );
  OAI22_X2 U11776 ( .A1(n6669), .A2(n11202), .B1(n12607), .B2(n11282), .ZN(
        pipeline_csr_N2163) );
  INV_X4 U11777 ( .A(pipeline_csr_N901), .ZN(n11203) );
  OAI22_X2 U11778 ( .A1(n6669), .A2(n11203), .B1(n12335), .B2(n11282), .ZN(
        pipeline_csr_N2162) );
  NAND2_X2 U11779 ( .A1(n9468), .A2(n12234), .ZN(n12244) );
  INV_X4 U11780 ( .A(pipeline_csr_N900), .ZN(n11204) );
  OAI22_X2 U11781 ( .A1(n12244), .A2(n11282), .B1(n6669), .B2(n11204), .ZN(
        pipeline_csr_N2161) );
  NAND2_X2 U11782 ( .A1(n9468), .A2(n12188), .ZN(n12196) );
  INV_X4 U11783 ( .A(pipeline_csr_N899), .ZN(n11205) );
  OAI22_X2 U11784 ( .A1(n12196), .A2(n11282), .B1(n6669), .B2(n11205), .ZN(
        pipeline_csr_N2160) );
  NAND2_X2 U11785 ( .A1(n9468), .A2(n12110), .ZN(n12118) );
  INV_X4 U11786 ( .A(pipeline_csr_N898), .ZN(n11206) );
  OAI22_X2 U11787 ( .A1(n12118), .A2(n11282), .B1(n6669), .B2(n11206), .ZN(
        pipeline_csr_N2159) );
  NAND2_X2 U11788 ( .A1(n9468), .A2(n12042), .ZN(n12050) );
  INV_X4 U11789 ( .A(pipeline_csr_N897), .ZN(n11207) );
  OAI22_X2 U11790 ( .A1(n12050), .A2(n11282), .B1(n6669), .B2(n11207), .ZN(
        pipeline_csr_N2158) );
  NAND2_X2 U11791 ( .A1(n9468), .A2(n11972), .ZN(n11980) );
  INV_X4 U11792 ( .A(pipeline_csr_N896), .ZN(n11208) );
  OAI22_X2 U11793 ( .A1(n11980), .A2(n11282), .B1(n6669), .B2(n11208), .ZN(
        pipeline_csr_N2157) );
  NAND2_X2 U11794 ( .A1(n9468), .A2(n11857), .ZN(n11865) );
  INV_X4 U11795 ( .A(pipeline_csr_N895), .ZN(n11209) );
  OAI22_X2 U11796 ( .A1(n11865), .A2(n11282), .B1(n6669), .B2(n11209), .ZN(
        pipeline_csr_N2156) );
  NAND2_X2 U11797 ( .A1(n9468), .A2(n11787), .ZN(n11797) );
  INV_X4 U11798 ( .A(pipeline_csr_N894), .ZN(n11210) );
  OAI22_X2 U11799 ( .A1(n11797), .A2(n11282), .B1(n6669), .B2(n11210), .ZN(
        pipeline_csr_N2155) );
  NAND2_X2 U11800 ( .A1(n9468), .A2(n11703), .ZN(n11713) );
  INV_X4 U11801 ( .A(pipeline_csr_N893), .ZN(n11211) );
  OAI22_X2 U11802 ( .A1(n11713), .A2(n11282), .B1(n6669), .B2(n11211), .ZN(
        pipeline_csr_N2154) );
  NAND2_X2 U11803 ( .A1(n9468), .A2(n11629), .ZN(n11639) );
  INV_X4 U11804 ( .A(pipeline_csr_N892), .ZN(n11212) );
  OAI22_X2 U11805 ( .A1(n11639), .A2(n11282), .B1(n6669), .B2(n11212), .ZN(
        pipeline_csr_N2153) );
  NAND2_X2 U11806 ( .A1(n9468), .A2(n11557), .ZN(n11567) );
  INV_X4 U11807 ( .A(pipeline_csr_N891), .ZN(n11213) );
  OAI22_X2 U11808 ( .A1(n11567), .A2(n11282), .B1(n6669), .B2(n11213), .ZN(
        pipeline_csr_N2152) );
  NAND2_X2 U11809 ( .A1(n9468), .A2(n11483), .ZN(n11493) );
  INV_X4 U11810 ( .A(pipeline_csr_N890), .ZN(n11214) );
  OAI22_X2 U11811 ( .A1(n11493), .A2(n11282), .B1(n6669), .B2(n11214), .ZN(
        pipeline_csr_N2151) );
  NAND2_X2 U11812 ( .A1(n9468), .A2(n11423), .ZN(n11433) );
  INV_X4 U11813 ( .A(pipeline_csr_N889), .ZN(n11215) );
  OAI22_X2 U11814 ( .A1(n11433), .A2(n11282), .B1(n6669), .B2(n11215), .ZN(
        pipeline_csr_N2150) );
  NAND2_X2 U11815 ( .A1(n9468), .A2(n11384), .ZN(n11394) );
  INV_X4 U11816 ( .A(pipeline_csr_N888), .ZN(n11216) );
  OAI22_X2 U11817 ( .A1(n11394), .A2(n11282), .B1(n6669), .B2(n11216), .ZN(
        pipeline_csr_N2149) );
  NAND2_X2 U11818 ( .A1(n9468), .A2(n11354), .ZN(n11364) );
  INV_X4 U11819 ( .A(pipeline_csr_N887), .ZN(n11217) );
  OAI22_X2 U11820 ( .A1(n11364), .A2(n11282), .B1(n6669), .B2(n11217), .ZN(
        pipeline_csr_N2148) );
  NAND2_X2 U11821 ( .A1(n9468), .A2(n11218), .ZN(n11330) );
  INV_X4 U11822 ( .A(pipeline_csr_N886), .ZN(n11219) );
  OAI22_X2 U11823 ( .A1(n11330), .A2(n11282), .B1(n6669), .B2(n11219), .ZN(
        pipeline_csr_N2147) );
  NAND2_X2 U11824 ( .A1(n9468), .A2(n11453), .ZN(n11463) );
  INV_X4 U11825 ( .A(pipeline_csr_N885), .ZN(n11220) );
  OAI22_X2 U11826 ( .A1(n11463), .A2(n11282), .B1(n6669), .B2(n11220), .ZN(
        pipeline_csr_N2146) );
  NAND2_X2 U11827 ( .A1(n9468), .A2(n11662), .ZN(n11672) );
  INV_X4 U11828 ( .A(pipeline_csr_N884), .ZN(n11221) );
  OAI22_X2 U11829 ( .A1(n11672), .A2(n11282), .B1(n6669), .B2(n11221), .ZN(
        pipeline_csr_N2145) );
  NAND2_X2 U11830 ( .A1(n9468), .A2(n11595), .ZN(n11605) );
  INV_X4 U11831 ( .A(pipeline_csr_N883), .ZN(n11222) );
  OAI22_X2 U11832 ( .A1(n11605), .A2(n11282), .B1(n6669), .B2(n11222), .ZN(
        pipeline_csr_N2144) );
  NAND2_X2 U11833 ( .A1(n9468), .A2(n11519), .ZN(n11529) );
  INV_X4 U11834 ( .A(pipeline_csr_N882), .ZN(n11223) );
  OAI22_X2 U11835 ( .A1(n11529), .A2(n11282), .B1(n6669), .B2(n11223), .ZN(
        pipeline_csr_N2143) );
  NAND2_X2 U11836 ( .A1(n9468), .A2(n12074), .ZN(n12084) );
  INV_X4 U11837 ( .A(pipeline_csr_N881), .ZN(n11224) );
  OAI22_X2 U11838 ( .A1(n12084), .A2(n11282), .B1(n6669), .B2(n11224), .ZN(
        pipeline_csr_N2142) );
  NAND2_X2 U11839 ( .A1(n9468), .A2(n11999), .ZN(n12009) );
  INV_X4 U11840 ( .A(pipeline_csr_N880), .ZN(n11225) );
  OAI22_X2 U11841 ( .A1(n12009), .A2(n11282), .B1(n6669), .B2(n11225), .ZN(
        pipeline_csr_N2141) );
  NAND2_X2 U11842 ( .A1(n9468), .A2(n11892), .ZN(n11941) );
  INV_X4 U11843 ( .A(pipeline_csr_N879), .ZN(n11226) );
  OAI22_X2 U11844 ( .A1(n11941), .A2(n11282), .B1(n6669), .B2(n11226), .ZN(
        pipeline_csr_N2140) );
  NAND2_X2 U11845 ( .A1(n9468), .A2(n11816), .ZN(n11826) );
  INV_X4 U11846 ( .A(pipeline_csr_N878), .ZN(n11227) );
  OAI22_X2 U11847 ( .A1(n11826), .A2(n11282), .B1(n6669), .B2(n11227), .ZN(
        pipeline_csr_N2139) );
  NAND2_X2 U11848 ( .A1(n9468), .A2(n11739), .ZN(n11754) );
  INV_X4 U11849 ( .A(pipeline_csr_N877), .ZN(n11228) );
  OAI22_X2 U11850 ( .A1(n11754), .A2(n11282), .B1(n6669), .B2(n11228), .ZN(
        pipeline_csr_N2138) );
  NAND2_X2 U11851 ( .A1(htif_pcr_req_data[4]), .A2(n13131), .ZN(n11252) );
  NAND2_X2 U11852 ( .A1(pipeline_regfile_N16), .A2(pipeline_dmem_type_2_), 
        .ZN(n11247) );
  NAND2_X2 U11853 ( .A1(pipeline_csr_mtvec[4]), .A2(n11229), .ZN(n11230) );
  OAI221_X2 U11854 ( .B1(n13105), .B2(n6836), .C1(n13098), .C2(n11231), .A(
        n11230), .ZN(n11232) );
  AOI221_X2 U11855 ( .B1(pipeline_csr_cycle_full[36]), .B2(n11233), .C1(
        pipeline_csr_time_full[4]), .C2(n6735), .A(n11232), .ZN(n11244) );
  AOI221_X2 U11857 ( .B1(pipeline_csr_instret_full[4]), .B2(n6640), .C1(n9527), 
        .C2(n11237), .A(n11236), .ZN(n11243) );
  OAI22_X2 U11858 ( .A1(n11264), .A2(n6827), .B1(n1487), .B2(n13114), .ZN(
        n11238) );
  AOI221_X2 U11859 ( .B1(pipeline_csr_cycle_full[4]), .B2(n13116), .C1(n11268), 
        .C2(n11239), .A(n11238), .ZN(n11242) );
  OAI22_X2 U11860 ( .A1(n13112), .A2(n12815), .B1(n1519), .B2(n9462), .ZN(
        n11240) );
  AOI221_X2 U11861 ( .B1(pipeline_csr_mtime_full[36]), .B2(n9528), .C1(n9466), 
        .C2(pipeline_csr_mtimecmp[4]), .A(n11240), .ZN(n11241) );
  NOR2_X2 U11862 ( .A1(n6713), .A2(n9463), .ZN(n11246) );
  NAND3_X2 U11863 ( .A1(n11247), .A2(n11246), .A3(n11245), .ZN(n11251) );
  NOR2_X2 U11864 ( .A1(n12522), .A2(n9467), .ZN(n11249) );
  NOR2_X2 U11865 ( .A1(n11280), .A2(n9270), .ZN(n11248) );
  NOR2_X2 U11866 ( .A1(n11249), .A2(n11248), .ZN(n11250) );
  NAND3_X2 U11867 ( .A1(n11252), .A2(n11251), .A3(n11250), .ZN(n12339) );
  NAND2_X2 U11868 ( .A1(n9468), .A2(n12339), .ZN(n12610) );
  INV_X4 U11869 ( .A(pipeline_csr_N876), .ZN(n11253) );
  OAI22_X2 U11870 ( .A1(n12610), .A2(n11282), .B1(n6669), .B2(n11253), .ZN(
        pipeline_csr_N2137) );
  INV_X4 U11871 ( .A(pipeline_csr_N875), .ZN(n11254) );
  OAI22_X2 U11872 ( .A1(n12147), .A2(n11282), .B1(n6669), .B2(n11254), .ZN(
        pipeline_csr_N2136) );
  INV_X4 U11873 ( .A(pipeline_csr_N874), .ZN(n11255) );
  OAI22_X2 U11874 ( .A1(n12260), .A2(n11282), .B1(n6669), .B2(n11255), .ZN(
        pipeline_csr_N2135) );
  INV_X4 U11875 ( .A(pipeline_csr_N873), .ZN(n11256) );
  OAI22_X2 U11876 ( .A1(n12354), .A2(n11282), .B1(n6669), .B2(n11256), .ZN(
        pipeline_csr_N2134) );
  NAND2_X2 U11877 ( .A1(pipeline_csr_time_full[32]), .A2(n11257), .ZN(n11258)
         );
  OAI221_X2 U11878 ( .B1(n13098), .B2(n11259), .C1(n13099), .C2(n6829), .A(
        n11258), .ZN(n11260) );
  AOI221_X2 U11879 ( .B1(pipeline_csr_time_full[0]), .B2(n6735), .C1(
        pipeline_csr_instret_full[0]), .C2(n6640), .A(n11260), .ZN(n11275) );
  OAI22_X2 U11880 ( .A1(n1447), .A2(n9464), .B1(n1255), .B2(n11261), .ZN(
        n11263) );
  AOI221_X2 U11881 ( .B1(pipeline_csr_from_host[0]), .B2(n9461), .C1(
        pipeline_csr_cycle_full[0]), .C2(n13116), .A(n11263), .ZN(n11274) );
  OAI22_X2 U11882 ( .A1(n11264), .A2(n6823), .B1(n1483), .B2(n13114), .ZN(
        n11265) );
  AOI221_X2 U11883 ( .B1(n11268), .B2(n11267), .C1(n11266), .C2(n12627), .A(
        n11265), .ZN(n11273) );
  INV_X4 U11884 ( .A(n13112), .ZN(n11741) );
  OAI22_X2 U11885 ( .A1(n1287), .A2(n11269), .B1(n13111), .B2(n6834), .ZN(
        n11270) );
  AOI221_X2 U11886 ( .B1(n6697), .B2(n11271), .C1(pipeline_csr_priv_stack_0), 
        .C2(n11741), .A(n11270), .ZN(n11272) );
  NAND4_X2 U11887 ( .A1(n11275), .A2(n11274), .A3(n11273), .A4(n11272), .ZN(
        n12630) );
  NAND2_X2 U11888 ( .A1(n6665), .A2(n12630), .ZN(n11276) );
  NAND2_X2 U11889 ( .A1(n9468), .A2(n12622), .ZN(n12614) );
  INV_X4 U11890 ( .A(pipeline_csr_N872), .ZN(n11281) );
  OAI22_X2 U11891 ( .A1(n12614), .A2(n11282), .B1(n6669), .B2(n11281), .ZN(
        pipeline_csr_N2133) );
  NOR2_X2 U11892 ( .A1(n11283), .A2(n11282), .ZN(n11285) );
  INV_X4 U11893 ( .A(pipeline_csr_N871), .ZN(n11286) );
  OAI22_X2 U11894 ( .A1(n6668), .A2(n11286), .B1(n12603), .B2(n11318), .ZN(
        pipeline_csr_N2132) );
  INV_X4 U11895 ( .A(pipeline_csr_N870), .ZN(n11287) );
  OAI22_X2 U11896 ( .A1(n6668), .A2(n11287), .B1(n12607), .B2(n11318), .ZN(
        pipeline_csr_N2131) );
  INV_X4 U11897 ( .A(pipeline_csr_N869), .ZN(n11288) );
  OAI22_X2 U11898 ( .A1(n6668), .A2(n11288), .B1(n12335), .B2(n11318), .ZN(
        pipeline_csr_N2130) );
  INV_X4 U11899 ( .A(pipeline_csr_N868), .ZN(n11289) );
  OAI22_X2 U11900 ( .A1(n12244), .A2(n11318), .B1(n6668), .B2(n11289), .ZN(
        pipeline_csr_N2129) );
  INV_X4 U11901 ( .A(pipeline_csr_N867), .ZN(n11290) );
  OAI22_X2 U11902 ( .A1(n12196), .A2(n11318), .B1(n6668), .B2(n11290), .ZN(
        pipeline_csr_N2128) );
  INV_X4 U11903 ( .A(pipeline_csr_N866), .ZN(n11291) );
  OAI22_X2 U11904 ( .A1(n12118), .A2(n11318), .B1(n6668), .B2(n11291), .ZN(
        pipeline_csr_N2127) );
  INV_X4 U11905 ( .A(pipeline_csr_N865), .ZN(n11292) );
  OAI22_X2 U11906 ( .A1(n12050), .A2(n11318), .B1(n6668), .B2(n11292), .ZN(
        pipeline_csr_N2126) );
  INV_X4 U11907 ( .A(pipeline_csr_N864), .ZN(n11293) );
  OAI22_X2 U11908 ( .A1(n11980), .A2(n11318), .B1(n6668), .B2(n11293), .ZN(
        pipeline_csr_N2125) );
  INV_X4 U11909 ( .A(pipeline_csr_N863), .ZN(n11294) );
  OAI22_X2 U11910 ( .A1(n11865), .A2(n11318), .B1(n6668), .B2(n11294), .ZN(
        pipeline_csr_N2124) );
  INV_X4 U11911 ( .A(pipeline_csr_N862), .ZN(n11295) );
  OAI22_X2 U11912 ( .A1(n6668), .A2(n11295), .B1(n11797), .B2(n11318), .ZN(
        pipeline_csr_N2123) );
  INV_X4 U11913 ( .A(pipeline_csr_N861), .ZN(n11296) );
  OAI22_X2 U11914 ( .A1(n11713), .A2(n11318), .B1(n6668), .B2(n11296), .ZN(
        pipeline_csr_N2122) );
  INV_X4 U11915 ( .A(pipeline_csr_N860), .ZN(n11297) );
  OAI22_X2 U11916 ( .A1(n11639), .A2(n11318), .B1(n6668), .B2(n11297), .ZN(
        pipeline_csr_N2121) );
  INV_X4 U11917 ( .A(pipeline_csr_N859), .ZN(n11298) );
  OAI22_X2 U11918 ( .A1(n11567), .A2(n11318), .B1(n6668), .B2(n11298), .ZN(
        pipeline_csr_N2120) );
  INV_X4 U11919 ( .A(pipeline_csr_N858), .ZN(n11299) );
  OAI22_X2 U11920 ( .A1(n11493), .A2(n11318), .B1(n6668), .B2(n11299), .ZN(
        pipeline_csr_N2119) );
  INV_X4 U11921 ( .A(pipeline_csr_N857), .ZN(n11300) );
  OAI22_X2 U11922 ( .A1(n11433), .A2(n11318), .B1(n6668), .B2(n11300), .ZN(
        pipeline_csr_N2118) );
  INV_X4 U11923 ( .A(pipeline_csr_N856), .ZN(n11301) );
  OAI22_X2 U11924 ( .A1(n11394), .A2(n11318), .B1(n6668), .B2(n11301), .ZN(
        pipeline_csr_N2117) );
  INV_X4 U11925 ( .A(pipeline_csr_N855), .ZN(n11302) );
  OAI22_X2 U11926 ( .A1(n11364), .A2(n11318), .B1(n6668), .B2(n11302), .ZN(
        pipeline_csr_N2116) );
  INV_X4 U11927 ( .A(pipeline_csr_N853), .ZN(n11303) );
  OAI22_X2 U11928 ( .A1(n11463), .A2(n11318), .B1(n6668), .B2(n11303), .ZN(
        pipeline_csr_N2114) );
  INV_X4 U11929 ( .A(pipeline_csr_N852), .ZN(n11304) );
  OAI22_X2 U11930 ( .A1(n11672), .A2(n11318), .B1(n6668), .B2(n11304), .ZN(
        pipeline_csr_N2113) );
  INV_X4 U11931 ( .A(pipeline_csr_N851), .ZN(n11305) );
  OAI22_X2 U11932 ( .A1(n11605), .A2(n11318), .B1(n6668), .B2(n11305), .ZN(
        pipeline_csr_N2112) );
  INV_X4 U11933 ( .A(pipeline_csr_N850), .ZN(n11306) );
  OAI22_X2 U11934 ( .A1(n11529), .A2(n11318), .B1(n6668), .B2(n11306), .ZN(
        pipeline_csr_N2111) );
  INV_X4 U11935 ( .A(pipeline_csr_N849), .ZN(n11307) );
  OAI22_X2 U11936 ( .A1(n12084), .A2(n11318), .B1(n6668), .B2(n11307), .ZN(
        pipeline_csr_N2110) );
  INV_X4 U11937 ( .A(pipeline_csr_N848), .ZN(n11308) );
  OAI22_X2 U11938 ( .A1(n12009), .A2(n11318), .B1(n6668), .B2(n11308), .ZN(
        pipeline_csr_N2109) );
  INV_X4 U11939 ( .A(pipeline_csr_N847), .ZN(n11309) );
  OAI22_X2 U11940 ( .A1(n11941), .A2(n11318), .B1(n6668), .B2(n11309), .ZN(
        pipeline_csr_N2108) );
  INV_X4 U11941 ( .A(pipeline_csr_N846), .ZN(n11310) );
  OAI22_X2 U11942 ( .A1(n11826), .A2(n11318), .B1(n6668), .B2(n11310), .ZN(
        pipeline_csr_N2107) );
  INV_X4 U11943 ( .A(pipeline_csr_N845), .ZN(n11311) );
  OAI22_X2 U11944 ( .A1(n11754), .A2(n11318), .B1(n6668), .B2(n11311), .ZN(
        pipeline_csr_N2106) );
  INV_X4 U11945 ( .A(pipeline_csr_N844), .ZN(n11312) );
  OAI22_X2 U11946 ( .A1(n12610), .A2(n11318), .B1(n6668), .B2(n11312), .ZN(
        pipeline_csr_N2105) );
  INV_X4 U11947 ( .A(pipeline_csr_N843), .ZN(n11313) );
  OAI22_X2 U11948 ( .A1(n12147), .A2(n11318), .B1(n6668), .B2(n11313), .ZN(
        pipeline_csr_N2104) );
  INV_X4 U11949 ( .A(pipeline_csr_N842), .ZN(n11314) );
  OAI22_X2 U11950 ( .A1(n12260), .A2(n11318), .B1(n6668), .B2(n11314), .ZN(
        pipeline_csr_N2103) );
  INV_X4 U11951 ( .A(pipeline_csr_N841), .ZN(n11315) );
  OAI22_X2 U11952 ( .A1(n12354), .A2(n11318), .B1(n6668), .B2(n11315), .ZN(
        pipeline_csr_N2102) );
  INV_X4 U11953 ( .A(pipeline_csr_N840), .ZN(n11316) );
  OAI22_X2 U11954 ( .A1(n12614), .A2(n11318), .B1(n6668), .B2(n11316), .ZN(
        pipeline_csr_N2101) );
  INV_X4 U11955 ( .A(pipeline_csr_N854), .ZN(n11317) );
  OAI22_X2 U11956 ( .A1(n11330), .A2(n11318), .B1(n6668), .B2(n11317), .ZN(
        pipeline_csr_N2115) );
  OAI22_X2 U11957 ( .A1(n6702), .A2(n11328), .B1(n11139), .B2(n9529), .ZN(
        n6162) );
  OAI22_X2 U11958 ( .A1(n6688), .A2(n11328), .B1(n1175), .B2(n3689), .ZN(n6130) );
  NAND3_X2 U11959 ( .A1(n6700), .A2(n9469), .A3(n6819), .ZN(n11319) );
  NAND2_X2 U11960 ( .A1(n9468), .A2(n11319), .ZN(n11321) );
  INV_X4 U11961 ( .A(pipeline_csr_N662), .ZN(n11322) );
  OAI22_X2 U11962 ( .A1(n12255), .A2(n11330), .B1(n6821), .B2(n11322), .ZN(
        pipeline_csr_N1902) );
  OAI22_X2 U11963 ( .A1(n6703), .A2(n11328), .B1(n11142), .B2(n3683), .ZN(
        n6067) );
  NAND2_X2 U11964 ( .A1(pipeline_csr_N822), .A2(n9476), .ZN(n11324) );
  OAI221_X2 U11965 ( .B1(n11328), .B2(n6704), .C1(n11143), .C2(n12352), .A(
        n11324), .ZN(n6000) );
  INV_X4 U11966 ( .A(pipeline_csr_N758), .ZN(n11325) );
  OAI22_X2 U11967 ( .A1(n9492), .A2(n11330), .B1(n9403), .B2(n11325), .ZN(
        pipeline_csr_N1998) );
  INV_X4 U11968 ( .A(pipeline_csr_N694), .ZN(n11326) );
  OAI22_X2 U11969 ( .A1(n9469), .A2(n11330), .B1(n9404), .B2(n11326), .ZN(
        pipeline_csr_N1934) );
  NAND2_X2 U11970 ( .A1(pipeline_csr_N790), .A2(n12346), .ZN(n11327) );
  OAI221_X2 U11971 ( .B1(n11328), .B2(n12347), .C1(n11145), .C2(n12349), .A(
        n11327), .ZN(n6032) );
  INV_X4 U11972 ( .A(pipeline_csr_N726), .ZN(n11329) );
  OAI22_X2 U11973 ( .A1(n12612), .A2(n11330), .B1(n9406), .B2(n11329), .ZN(
        pipeline_csr_N1966) );
  OAI22_X2 U11974 ( .A1(n7197), .A2(n6691), .B1(n436), .B2(n9525), .ZN(n6348)
         );
  NAND2_X2 U11975 ( .A1(n9471), .A2(pipeline_alu_src_a[24]), .ZN(n12032) );
  NAND2_X2 U11976 ( .A1(n12276), .A2(n6608), .ZN(n12177) );
  NAND2_X2 U11977 ( .A1(n11869), .A2(n6560), .ZN(n12307) );
  NAND2_X2 U11978 ( .A1(n9489), .A2(n6980), .ZN(n11843) );
  NAND4_X2 U11979 ( .A1(n12032), .A2(n12177), .A3(n12307), .A4(n11843), .ZN(
        n11576) );
  NAND2_X2 U11980 ( .A1(n9471), .A2(n6565), .ZN(n12309) );
  NAND2_X2 U11981 ( .A1(n12276), .A2(pipeline_alu_src_a[29]), .ZN(n12571) );
  NAND2_X2 U11982 ( .A1(n11869), .A2(n6997), .ZN(n11331) );
  NAND4_X2 U11983 ( .A1(n12309), .A2(n12571), .A3(n11331), .A4(n12175), .ZN(
        n11577) );
  NAND2_X2 U11984 ( .A1(n11869), .A2(pipeline_alu_src_a[18]), .ZN(n11690) );
  INV_X4 U11985 ( .A(n11877), .ZN(n12133) );
  NAND2_X2 U11986 ( .A1(n9471), .A2(pipeline_alu_src_a[20]), .ZN(n11692) );
  NAND2_X2 U11987 ( .A1(n12276), .A2(pipeline_alu_src_a[21]), .ZN(n11845) );
  NAND2_X2 U11988 ( .A1(n9489), .A2(pipeline_alu_src_a[19]), .ZN(n11333) );
  NAND2_X2 U11989 ( .A1(n11869), .A2(n6625), .ZN(n12030) );
  NAND4_X2 U11990 ( .A1(n11692), .A2(n11845), .A3(n11333), .A4(n12030), .ZN(
        n11876) );
  INV_X4 U11991 ( .A(n11876), .ZN(n11543) );
  OAI22_X2 U11992 ( .A1(n12133), .A2(n9509), .B1(n11543), .B2(n9507), .ZN(
        n11334) );
  AOI221_X2 U11993 ( .B1(n9511), .B2(n11576), .C1(n12780), .C2(n11577), .A(
        n11334), .ZN(n11335) );
  NAND2_X2 U11994 ( .A1(n9489), .A2(n7005), .ZN(n11834) );
  OAI22_X2 U11995 ( .A1(n11335), .A2(n12772), .B1(n11834), .B2(n11645), .ZN(
        n11340) );
  INV_X4 U11996 ( .A(n12659), .ZN(n11339) );
  NOR2_X2 U11997 ( .A1(pipeline_alu_src_b[15]), .A2(n12357), .ZN(n11336) );
  NOR2_X2 U11998 ( .A1(n9513), .A2(n11336), .ZN(n11337) );
  NOR2_X2 U11999 ( .A1(n11414), .A2(n11337), .ZN(n11338) );
  NOR3_X2 U12000 ( .A1(n11340), .A2(n11339), .A3(n11338), .ZN(n11351) );
  NAND4_X2 U12001 ( .A1(n12131), .A2(n11717), .A3(n11870), .A4(n12367), .ZN(
        n11827) );
  INV_X4 U12002 ( .A(n11827), .ZN(n11532) );
  NAND2_X2 U12003 ( .A1(n12276), .A2(n6632), .ZN(n11342) );
  NAND2_X2 U12004 ( .A1(n9489), .A2(n6634), .ZN(n12129) );
  NAND4_X2 U12005 ( .A1(n11342), .A2(n12369), .A3(n12129), .A4(n11341), .ZN(
        n12126) );
  INV_X4 U12006 ( .A(n12126), .ZN(n11535) );
  AOI221_X2 U12007 ( .B1(n9471), .B2(n11570), .C1(n12276), .C2(n11573), .A(
        n11343), .ZN(n11830) );
  NAND2_X2 U12008 ( .A1(n12276), .A2(n6972), .ZN(n11872) );
  NAND4_X2 U12009 ( .A1(n11872), .A2(n11721), .A3(n11569), .A4(n11715), .ZN(
        n11829) );
  OAI22_X2 U12010 ( .A1(n11830), .A2(n9509), .B1(n9507), .B2(n11829), .ZN(
        n11344) );
  AOI221_X2 U12011 ( .B1(n11532), .B2(n9511), .C1(n11535), .C2(n12780), .A(
        n11344), .ZN(n12584) );
  INV_X4 U12012 ( .A(n12584), .ZN(n11348) );
  MUX2_X2 U12013 ( .A(n12793), .B(n9479), .S(n11414), .Z(n11345) );
  NOR2_X2 U12014 ( .A1(n9513), .A2(n11345), .ZN(n11346) );
  OAI22_X2 U12015 ( .A1(n12785), .A2(n11348), .B1(n11347), .B2(n11346), .ZN(
        n11349) );
  AOI221_X2 U12016 ( .B1(pipeline_alu_N74), .B2(n6813), .C1(pipeline_alu_N268), 
        .C2(n6812), .A(n11349), .ZN(n11350) );
  NAND2_X2 U12017 ( .A1(n11351), .A2(n11350), .ZN(dmem_haddr[15]) );
  MUX2_X2 U12018 ( .A(pipeline_alu_out_WB[15]), .B(dmem_haddr[15]), .S(n9523), 
        .Z(n5829) );
  OAI22_X2 U12019 ( .A1(n9515), .A2(n11352), .B1(n550), .B2(n9498), .ZN(n11353) );
  AOI221_X2 U12020 ( .B1(n12668), .B2(n11354), .C1(pipeline_alu_out_WB[15]), 
        .C2(n12809), .A(n11353), .ZN(n11355) );
  INV_X4 U12021 ( .A(n11355), .ZN(n5797) );
  NAND2_X2 U12022 ( .A1(pipeline_csr_N316), .A2(n6750), .ZN(n11356) );
  OAI221_X2 U12023 ( .B1(n11362), .B2(n6705), .C1(n1498), .C2(n6687), .A(
        n11356), .ZN(n5860) );
  OAI22_X2 U12024 ( .A1(n6659), .A2(n11362), .B1(n1270), .B2(n6689), .ZN(n6096) );
  OAI22_X2 U12025 ( .A1(n6703), .A2(n11362), .B1(n1238), .B2(n3683), .ZN(n6066) );
  INV_X4 U12026 ( .A(pipeline_csr_N759), .ZN(n11357) );
  OAI22_X2 U12027 ( .A1(n9492), .A2(n11364), .B1(n9403), .B2(n11357), .ZN(
        pipeline_csr_N1999) );
  NAND2_X2 U12028 ( .A1(pipeline_csr_N823), .A2(n9476), .ZN(n11358) );
  OAI221_X2 U12029 ( .B1(n11362), .B2(n6704), .C1(n1430), .C2(n12352), .A(
        n11358), .ZN(n5999) );
  OAI22_X2 U12030 ( .A1(n6702), .A2(n11362), .B1(n11107), .B2(n9529), .ZN(
        n6161) );
  OAI22_X2 U12031 ( .A1(n6688), .A2(n11362), .B1(n1176), .B2(n9530), .ZN(n6129) );
  INV_X4 U12032 ( .A(pipeline_csr_N727), .ZN(n11359) );
  OAI22_X2 U12033 ( .A1(n12612), .A2(n11364), .B1(n9405), .B2(n11359), .ZN(
        pipeline_csr_N1967) );
  INV_X4 U12034 ( .A(pipeline_csr_N663), .ZN(n11360) );
  OAI22_X2 U12035 ( .A1(n12255), .A2(n11364), .B1(n6821), .B2(n11360), .ZN(
        pipeline_csr_N1903) );
  NAND2_X2 U12036 ( .A1(pipeline_csr_N791), .A2(n12346), .ZN(n11361) );
  OAI221_X2 U12037 ( .B1(n11362), .B2(n12347), .C1(n11109), .C2(n12349), .A(
        n11361), .ZN(n6031) );
  INV_X4 U12038 ( .A(pipeline_csr_N695), .ZN(n11363) );
  OAI22_X2 U12039 ( .A1(n9469), .A2(n11364), .B1(n9404), .B2(n11363), .ZN(
        pipeline_csr_N1935) );
  OAI22_X2 U12040 ( .A1(n7189), .A2(n6691), .B1(n438), .B2(n9523), .ZN(n6349)
         );
  INV_X4 U12041 ( .A(n11366), .ZN(n11944) );
  AOI221_X2 U12042 ( .B1(n9471), .B2(n6613), .C1(n12276), .C2(n11510), .A(
        n11367), .ZN(n11653) );
  INV_X4 U12043 ( .A(n11653), .ZN(n11950) );
  NAND2_X2 U12044 ( .A1(n11946), .A2(n9511), .ZN(n11369) );
  MUX2_X2 U12045 ( .A(n12355), .B(n12357), .S(n11474), .Z(n11370) );
  NAND2_X2 U12046 ( .A1(n11370), .A2(n9512), .ZN(n11375) );
  NOR2_X2 U12047 ( .A1(n9513), .A2(n11371), .ZN(n11373) );
  NAND2_X2 U12048 ( .A1(n12662), .A2(pipeline_alu_src_b[4]), .ZN(n11407) );
  AOI221_X2 U12049 ( .B1(n9471), .B2(n11414), .C1(n12276), .C2(n11570), .A(
        n11377), .ZN(n11947) );
  INV_X4 U12050 ( .A(n11947), .ZN(n12221) );
  OAI22_X2 U12051 ( .A1(n11378), .A2(n12772), .B1(n12182), .B2(n12221), .ZN(
        n11379) );
  AOI221_X2 U12052 ( .B1(pipeline_alu_N75), .B2(n6813), .C1(pipeline_alu_N269), 
        .C2(n6812), .A(n11379), .ZN(n11380) );
  NAND2_X2 U12053 ( .A1(n11381), .A2(n11380), .ZN(dmem_haddr[16]) );
  MUX2_X2 U12054 ( .A(pipeline_alu_out_WB[16]), .B(dmem_haddr[16]), .S(n9524), 
        .Z(n5828) );
  OAI22_X2 U12055 ( .A1(n9515), .A2(n11382), .B1(n551), .B2(n9498), .ZN(n11383) );
  AOI221_X2 U12056 ( .B1(n12668), .B2(n11384), .C1(pipeline_alu_out_WB[16]), 
        .C2(n12809), .A(n11383), .ZN(n11385) );
  INV_X4 U12057 ( .A(n11385), .ZN(n5796) );
  NAND2_X2 U12058 ( .A1(pipeline_csr_N317), .A2(n6750), .ZN(n11386) );
  OAI221_X2 U12059 ( .B1(n11392), .B2(n6705), .C1(n1499), .C2(n6687), .A(
        n11386), .ZN(n5859) );
  OAI22_X2 U12060 ( .A1(n6659), .A2(n11392), .B1(n1271), .B2(n6689), .ZN(n6097) );
  OAI22_X2 U12061 ( .A1(n6702), .A2(n11392), .B1(n11081), .B2(n9529), .ZN(
        n6160) );
  OAI22_X2 U12062 ( .A1(n6688), .A2(n11392), .B1(n1177), .B2(n9530), .ZN(n6128) );
  INV_X4 U12063 ( .A(pipeline_csr_N664), .ZN(n11387) );
  OAI22_X2 U12064 ( .A1(n12255), .A2(n11394), .B1(n6821), .B2(n11387), .ZN(
        pipeline_csr_N1904) );
  OAI22_X2 U12065 ( .A1(n6703), .A2(n11392), .B1(n11084), .B2(n3683), .ZN(
        n6065) );
  NAND2_X2 U12066 ( .A1(pipeline_csr_N824), .A2(n9476), .ZN(n11388) );
  OAI221_X2 U12067 ( .B1(n11392), .B2(n6704), .C1(n11085), .C2(n12352), .A(
        n11388), .ZN(n5998) );
  INV_X4 U12068 ( .A(pipeline_csr_N760), .ZN(n11389) );
  OAI22_X2 U12069 ( .A1(n9492), .A2(n11394), .B1(n9403), .B2(n11389), .ZN(
        pipeline_csr_N2000) );
  INV_X4 U12070 ( .A(pipeline_csr_N696), .ZN(n11390) );
  OAI22_X2 U12071 ( .A1(n9469), .A2(n11394), .B1(n12257), .B2(n11390), .ZN(
        pipeline_csr_N1936) );
  NAND2_X2 U12072 ( .A1(pipeline_csr_N792), .A2(n12346), .ZN(n11391) );
  OAI221_X2 U12073 ( .B1(n11392), .B2(n12347), .C1(n11087), .C2(n12349), .A(
        n11391), .ZN(n6030) );
  INV_X4 U12074 ( .A(pipeline_csr_N728), .ZN(n11393) );
  OAI22_X2 U12075 ( .A1(n12612), .A2(n11394), .B1(n9405), .B2(n11393), .ZN(
        pipeline_csr_N1968) );
  OAI22_X2 U12076 ( .A1(n7196), .A2(n6691), .B1(n440), .B2(n9524), .ZN(n6350)
         );
  NAND2_X2 U12077 ( .A1(n12199), .A2(n12800), .ZN(n12089) );
  INV_X4 U12078 ( .A(n12089), .ZN(n12165) );
  NAND2_X2 U12079 ( .A1(n9471), .A2(n6561), .ZN(n12178) );
  NAND2_X2 U12080 ( .A1(n9489), .A2(n6609), .ZN(n12029) );
  NAND2_X2 U12081 ( .A1(n11869), .A2(n6564), .ZN(n12570) );
  NAND4_X2 U12082 ( .A1(n12308), .A2(n12178), .A3(n12029), .A4(n12570), .ZN(
        n12019) );
  INV_X4 U12083 ( .A(n12019), .ZN(n11680) );
  NOR2_X2 U12084 ( .A1(pipeline_alu_src_a[29]), .A2(n12565), .ZN(n11395) );
  NOR2_X2 U12085 ( .A1(n11869), .A2(n11395), .ZN(n11396) );
  NAND2_X2 U12086 ( .A1(n12276), .A2(pipeline_alu_src_a[19]), .ZN(n11691) );
  NAND2_X2 U12087 ( .A1(n9471), .A2(pipeline_alu_src_a[18]), .ZN(n11398) );
  NAND2_X2 U12088 ( .A1(n11869), .A2(pipeline_alu_src_a[20]), .ZN(n11844) );
  NAND4_X2 U12089 ( .A1(n11691), .A2(n11398), .A3(n11397), .A4(n11844), .ZN(
        n12057) );
  NAND2_X2 U12090 ( .A1(n12276), .A2(n6980), .ZN(n12031) );
  NAND2_X2 U12091 ( .A1(n9471), .A2(n6625), .ZN(n11846) );
  NAND2_X2 U12092 ( .A1(n9489), .A2(pipeline_alu_src_a[21]), .ZN(n11689) );
  NAND2_X2 U12093 ( .A1(n11869), .A2(pipeline_alu_src_a[24]), .ZN(n12176) );
  NAND4_X2 U12094 ( .A1(n12031), .A2(n11846), .A3(n11689), .A4(n12176), .ZN(
        n12056) );
  OAI22_X2 U12095 ( .A1(n9509), .A2(n12057), .B1(n9507), .B2(n12056), .ZN(
        n11399) );
  AOI221_X2 U12096 ( .B1(n11680), .B2(n9511), .C1(n12780), .C2(n11679), .A(
        n11399), .ZN(n12364) );
  NAND2_X2 U12097 ( .A1(n12276), .A2(n6635), .ZN(n12370) );
  NAND4_X2 U12098 ( .A1(n12132), .A2(n12370), .A3(n11400), .A4(n11716), .ZN(
        n12013) );
  INV_X4 U12099 ( .A(n12013), .ZN(n11443) );
  INV_X4 U12100 ( .A(n11675), .ZN(n12017) );
  NAND4_X2 U12101 ( .A1(n11873), .A2(n11718), .A3(n12130), .A4(n11719), .ZN(
        n12010) );
  NAND2_X2 U12102 ( .A1(n9511), .A2(n12010), .ZN(n11402) );
  NOR2_X2 U12103 ( .A1(pipeline_alu_src_b[17]), .A2(n12357), .ZN(n11403) );
  NOR2_X2 U12104 ( .A1(n9513), .A2(n11403), .ZN(n11408) );
  NAND2_X2 U12105 ( .A1(n11406), .A2(n11405), .ZN(n11673) );
  INV_X4 U12106 ( .A(n11407), .ZN(n12174) );
  NAND2_X2 U12107 ( .A1(n12174), .A2(n9510), .ZN(n11534) );
  OAI221_X2 U12108 ( .B1(n11546), .B2(n11408), .C1(n11673), .C2(n11534), .A(
        n12659), .ZN(n11409) );
  AOI221_X2 U12109 ( .B1(n12165), .B2(n12364), .C1(n12172), .C2(n11410), .A(
        n11409), .ZN(n11420) );
  NAND2_X2 U12110 ( .A1(n9489), .A2(pipeline_alu_src_a[29]), .ZN(n12306) );
  NAND2_X2 U12111 ( .A1(n9471), .A2(n6997), .ZN(n12572) );
  NAND3_X2 U12112 ( .A1(n12306), .A2(n12572), .A3(n11411), .ZN(n12025) );
  INV_X4 U12113 ( .A(n12057), .ZN(n11437) );
  INV_X4 U12114 ( .A(n12056), .ZN(n11681) );
  OAI22_X2 U12115 ( .A1(n11437), .A2(n9509), .B1(n11681), .B2(n9507), .ZN(
        n11412) );
  AOI221_X2 U12116 ( .B1(n9511), .B2(n12019), .C1(n12780), .C2(n12025), .A(
        n11412), .ZN(n12366) );
  INV_X4 U12117 ( .A(n12014), .ZN(n12317) );
  MUX2_X2 U12118 ( .A(n12355), .B(n12357), .S(n11546), .Z(n11415) );
  NAND2_X2 U12119 ( .A1(n11415), .A2(n9512), .ZN(n11416) );
  NAND2_X2 U12120 ( .A1(n11416), .A2(pipeline_alu_src_b[17]), .ZN(n11417) );
  OAI221_X2 U12121 ( .B1(n12366), .B2(n12639), .C1(n12182), .C2(n12317), .A(
        n11417), .ZN(n11418) );
  AOI221_X2 U12122 ( .B1(pipeline_alu_N76), .B2(n6813), .C1(pipeline_alu_N270), 
        .C2(n6812), .A(n11418), .ZN(n11419) );
  NAND2_X2 U12123 ( .A1(n11420), .A2(n11419), .ZN(dmem_haddr[17]) );
  MUX2_X2 U12124 ( .A(pipeline_alu_out_WB[17]), .B(dmem_haddr[17]), .S(n9524), 
        .Z(n5827) );
  OAI22_X2 U12125 ( .A1(n12805), .A2(n11421), .B1(n552), .B2(n9498), .ZN(
        n11422) );
  AOI221_X2 U12126 ( .B1(n12668), .B2(n11423), .C1(pipeline_alu_out_WB[17]), 
        .C2(n12809), .A(n11422), .ZN(n11424) );
  INV_X4 U12127 ( .A(n11424), .ZN(n5795) );
  NAND2_X2 U12128 ( .A1(pipeline_csr_N318), .A2(n6750), .ZN(n11425) );
  OAI221_X2 U12129 ( .B1(n11431), .B2(n6705), .C1(n1500), .C2(n6687), .A(
        n11425), .ZN(n5858) );
  OAI22_X2 U12130 ( .A1(n6659), .A2(n11431), .B1(n1272), .B2(n6689), .ZN(n6098) );
  OAI22_X2 U12131 ( .A1(n6702), .A2(n11431), .B1(n11054), .B2(n9529), .ZN(
        n6159) );
  OAI22_X2 U12132 ( .A1(n6688), .A2(n11431), .B1(n1178), .B2(n3689), .ZN(n6127) );
  INV_X4 U12133 ( .A(pipeline_csr_N665), .ZN(n11426) );
  OAI22_X2 U12134 ( .A1(n12255), .A2(n11433), .B1(n6821), .B2(n11426), .ZN(
        pipeline_csr_N1905) );
  OAI22_X2 U12135 ( .A1(n6703), .A2(n11431), .B1(n11057), .B2(n3683), .ZN(
        n6064) );
  NAND2_X2 U12136 ( .A1(pipeline_csr_N825), .A2(n9476), .ZN(n11427) );
  OAI221_X2 U12137 ( .B1(n11431), .B2(n6704), .C1(n11058), .C2(n12352), .A(
        n11427), .ZN(n5997) );
  INV_X4 U12138 ( .A(pipeline_csr_N761), .ZN(n11428) );
  OAI22_X2 U12139 ( .A1(n9492), .A2(n11433), .B1(n9403), .B2(n11428), .ZN(
        pipeline_csr_N2001) );
  INV_X4 U12140 ( .A(pipeline_csr_N697), .ZN(n11429) );
  OAI22_X2 U12141 ( .A1(n9469), .A2(n11433), .B1(n9404), .B2(n11429), .ZN(
        pipeline_csr_N1937) );
  NAND2_X2 U12142 ( .A1(pipeline_csr_N793), .A2(n12346), .ZN(n11430) );
  OAI221_X2 U12143 ( .B1(n11431), .B2(n12347), .C1(n11060), .C2(n12349), .A(
        n11430), .ZN(n6029) );
  INV_X4 U12144 ( .A(pipeline_csr_N729), .ZN(n11432) );
  OAI22_X2 U12145 ( .A1(n12612), .A2(n11433), .B1(n9406), .B2(n11432), .ZN(
        pipeline_csr_N1969) );
  OAI22_X2 U12146 ( .A1(n7195), .A2(n6691), .B1(n442), .B2(n9525), .ZN(n6351)
         );
  NAND2_X2 U12147 ( .A1(n9479), .A2(n11446), .ZN(n11434) );
  NAND2_X2 U12148 ( .A1(n11434), .A2(n9512), .ZN(n11441) );
  NAND2_X2 U12149 ( .A1(n9510), .A2(n12025), .ZN(n11435) );
  NAND2_X2 U12150 ( .A1(n11435), .A2(n11641), .ZN(n12322) );
  OAI22_X2 U12151 ( .A1(n12371), .A2(n12776), .B1(n11437), .B2(n9507), .ZN(
        n11438) );
  AOI221_X2 U12152 ( .B1(n9511), .B2(n12056), .C1(n12780), .C2(n12019), .A(
        n11438), .ZN(n11439) );
  OAI22_X2 U12153 ( .A1(n11439), .A2(n12772), .B1(n11679), .B2(n11645), .ZN(
        n11440) );
  AOI221_X2 U12154 ( .B1(n11441), .B2(n6568), .C1(n12062), .C2(n12322), .A(
        n11440), .ZN(n11450) );
  OAI22_X2 U12155 ( .A1(n11675), .A2(n9509), .B1(n9507), .B2(n12010), .ZN(
        n11442) );
  AOI221_X2 U12156 ( .B1(n11443), .B2(n9511), .C1(n12780), .C2(n11673), .A(
        n11442), .ZN(n12319) );
  INV_X4 U12157 ( .A(n12319), .ZN(n11447) );
  MUX2_X2 U12158 ( .A(n12793), .B(n9479), .S(n11573), .Z(n11444) );
  NOR2_X2 U12159 ( .A1(n9513), .A2(n11444), .ZN(n11445) );
  OAI22_X2 U12160 ( .A1(n12785), .A2(n11447), .B1(n11446), .B2(n11445), .ZN(
        n11448) );
  AOI221_X2 U12161 ( .B1(pipeline_alu_N72), .B2(n6813), .C1(pipeline_alu_N266), 
        .C2(n6812), .A(n11448), .ZN(n11449) );
  NAND2_X2 U12162 ( .A1(n11450), .A2(n11449), .ZN(dmem_haddr[13]) );
  MUX2_X2 U12163 ( .A(pipeline_alu_out_WB[13]), .B(dmem_haddr[13]), .S(n9522), 
        .Z(n5831) );
  OAI22_X2 U12164 ( .A1(n12805), .A2(n11451), .B1(n548), .B2(n9498), .ZN(
        n11452) );
  AOI221_X2 U12165 ( .B1(n12668), .B2(n11453), .C1(pipeline_alu_out_WB[13]), 
        .C2(n12809), .A(n11452), .ZN(n11454) );
  INV_X4 U12166 ( .A(n11454), .ZN(n5799) );
  NAND2_X2 U12167 ( .A1(pipeline_csr_N314), .A2(n6750), .ZN(n11455) );
  OAI221_X2 U12168 ( .B1(n11461), .B2(n6705), .C1(n1496), .C2(n6687), .A(
        n11455), .ZN(n5862) );
  OAI22_X2 U12169 ( .A1(n6659), .A2(n11461), .B1(n1268), .B2(n6689), .ZN(n6094) );
  OAI22_X2 U12170 ( .A1(n6702), .A2(n11461), .B1(n11027), .B2(n9529), .ZN(
        n6163) );
  OAI22_X2 U12171 ( .A1(n6688), .A2(n11461), .B1(n1174), .B2(n3689), .ZN(n6131) );
  INV_X4 U12172 ( .A(pipeline_csr_N661), .ZN(n11456) );
  OAI22_X2 U12173 ( .A1(n12255), .A2(n11463), .B1(n6821), .B2(n11456), .ZN(
        pipeline_csr_N1901) );
  OAI22_X2 U12174 ( .A1(n6703), .A2(n11461), .B1(n11030), .B2(n3683), .ZN(
        n6068) );
  NAND2_X2 U12175 ( .A1(pipeline_csr_N821), .A2(n9476), .ZN(n11457) );
  OAI221_X2 U12176 ( .B1(n11461), .B2(n6704), .C1(n11031), .C2(n12352), .A(
        n11457), .ZN(n6001) );
  INV_X4 U12177 ( .A(pipeline_csr_N757), .ZN(n11458) );
  OAI22_X2 U12178 ( .A1(n9492), .A2(n11463), .B1(n9403), .B2(n11458), .ZN(
        pipeline_csr_N1997) );
  INV_X4 U12179 ( .A(pipeline_csr_N693), .ZN(n11459) );
  OAI22_X2 U12180 ( .A1(n9469), .A2(n11463), .B1(n12257), .B2(n11459), .ZN(
        pipeline_csr_N1933) );
  NAND2_X2 U12181 ( .A1(pipeline_csr_N789), .A2(n12346), .ZN(n11460) );
  OAI221_X2 U12182 ( .B1(n11461), .B2(n12347), .C1(n11033), .C2(n12349), .A(
        n11460), .ZN(n6033) );
  INV_X4 U12183 ( .A(pipeline_csr_N725), .ZN(n11462) );
  OAI22_X2 U12184 ( .A1(n12612), .A2(n11463), .B1(n9406), .B2(n11462), .ZN(
        pipeline_csr_N1965) );
  OAI22_X2 U12185 ( .A1(n7198), .A2(n6691), .B1(n434), .B2(n9523), .ZN(n6347)
         );
  INV_X4 U12186 ( .A(n11495), .ZN(n11763) );
  OAI22_X2 U12187 ( .A1(n12776), .A2(n11801), .B1(n9507), .B2(n11500), .ZN(
        n11464) );
  AOI221_X2 U12188 ( .B1(n11763), .B2(n9511), .C1(n12780), .C2(n11501), .A(
        n11464), .ZN(n12269) );
  INV_X4 U12189 ( .A(n11758), .ZN(n12087) );
  NAND2_X2 U12190 ( .A1(n11757), .A2(n9511), .ZN(n11465) );
  NOR2_X2 U12191 ( .A1(pipeline_alu_src_b[18]), .A2(n12357), .ZN(n11467) );
  NOR2_X2 U12192 ( .A1(n9513), .A2(n11467), .ZN(n11468) );
  OAI221_X2 U12193 ( .B1(n11547), .B2(n11468), .C1(n11507), .C2(n11534), .A(
        n12659), .ZN(n11469) );
  AOI221_X2 U12194 ( .B1(n12165), .B2(n12269), .C1(n12172), .C2(n11470), .A(
        n11469), .ZN(n11480) );
  INV_X4 U12195 ( .A(n11500), .ZN(n11764) );
  OAI22_X2 U12196 ( .A1(n11471), .A2(n9509), .B1(n11764), .B2(n9507), .ZN(
        n11472) );
  AOI221_X2 U12197 ( .B1(n9511), .B2(n11495), .C1(n12780), .C2(n11770), .A(
        n11472), .ZN(n12271) );
  INV_X4 U12198 ( .A(n12647), .ZN(n11760) );
  MUX2_X2 U12199 ( .A(n12355), .B(n12357), .S(n11547), .Z(n11475) );
  NAND2_X2 U12200 ( .A1(n11475), .A2(n9512), .ZN(n11476) );
  NAND2_X2 U12201 ( .A1(n11476), .A2(pipeline_alu_src_b[18]), .ZN(n11477) );
  OAI221_X2 U12202 ( .B1(n12271), .B2(n12639), .C1(n11760), .C2(n12182), .A(
        n11477), .ZN(n11478) );
  AOI221_X2 U12203 ( .B1(pipeline_alu_N77), .B2(n6813), .C1(pipeline_alu_N271), 
        .C2(n6812), .A(n11478), .ZN(n11479) );
  NAND2_X2 U12204 ( .A1(n11480), .A2(n11479), .ZN(dmem_haddr[18]) );
  MUX2_X2 U12205 ( .A(pipeline_alu_out_WB[18]), .B(dmem_haddr[18]), .S(n9524), 
        .Z(n5826) );
  OAI22_X2 U12206 ( .A1(n12805), .A2(n11481), .B1(n553), .B2(n9498), .ZN(
        n11482) );
  AOI221_X2 U12207 ( .B1(n12668), .B2(n11483), .C1(pipeline_alu_out_WB[18]), 
        .C2(n12809), .A(n11482), .ZN(n11484) );
  INV_X4 U12208 ( .A(n11484), .ZN(n5794) );
  NAND2_X2 U12209 ( .A1(pipeline_csr_N319), .A2(n6750), .ZN(n11485) );
  OAI221_X2 U12210 ( .B1(n11491), .B2(n6705), .C1(n1501), .C2(n6687), .A(
        n11485), .ZN(n5857) );
  OAI22_X2 U12211 ( .A1(n6659), .A2(n11491), .B1(n1273), .B2(n6689), .ZN(n6099) );
  OAI22_X2 U12212 ( .A1(n6702), .A2(n11491), .B1(n11005), .B2(n9529), .ZN(
        n6158) );
  OAI22_X2 U12213 ( .A1(n6688), .A2(n11491), .B1(n1179), .B2(n3689), .ZN(n6126) );
  INV_X4 U12214 ( .A(pipeline_csr_N666), .ZN(n11486) );
  OAI22_X2 U12215 ( .A1(n12255), .A2(n11493), .B1(n6821), .B2(n11486), .ZN(
        pipeline_csr_N1906) );
  OAI22_X2 U12216 ( .A1(n6703), .A2(n11491), .B1(n10997), .B2(n3683), .ZN(
        n6063) );
  NAND2_X2 U12217 ( .A1(pipeline_csr_N826), .A2(n9476), .ZN(n11487) );
  OAI221_X2 U12218 ( .B1(n11491), .B2(n6704), .C1(n10998), .C2(n12352), .A(
        n11487), .ZN(n5996) );
  INV_X4 U12219 ( .A(pipeline_csr_N762), .ZN(n11488) );
  OAI22_X2 U12220 ( .A1(n9492), .A2(n11493), .B1(n9403), .B2(n11488), .ZN(
        pipeline_csr_N2002) );
  INV_X4 U12221 ( .A(pipeline_csr_N698), .ZN(n11489) );
  OAI22_X2 U12222 ( .A1(n9469), .A2(n11493), .B1(n12257), .B2(n11489), .ZN(
        pipeline_csr_N1938) );
  NAND2_X2 U12223 ( .A1(pipeline_csr_N794), .A2(n12346), .ZN(n11490) );
  OAI221_X2 U12224 ( .B1(n11491), .B2(n12347), .C1(n11000), .C2(n12349), .A(
        n11490), .ZN(n6028) );
  INV_X4 U12225 ( .A(pipeline_csr_N730), .ZN(n11492) );
  OAI22_X2 U12226 ( .A1(n12612), .A2(n11493), .B1(n9405), .B2(n11492), .ZN(
        pipeline_csr_N1970) );
  OAI22_X2 U12227 ( .A1(n7188), .A2(n6691), .B1(n444), .B2(n9525), .ZN(n6352)
         );
  NAND2_X2 U12228 ( .A1(n9479), .A2(n11513), .ZN(n11494) );
  NAND2_X2 U12229 ( .A1(n11494), .A2(n9512), .ZN(n11506) );
  NAND2_X2 U12230 ( .A1(n9508), .A2(n11770), .ZN(n11496) );
  NAND2_X2 U12231 ( .A1(n9510), .A2(n11495), .ZN(n11502) );
  NAND3_X2 U12232 ( .A1(n11496), .A2(n11502), .A3(n12027), .ZN(n12094) );
  OAI22_X2 U12233 ( .A1(n11510), .A2(n12565), .B1(n11573), .B2(n9400), .ZN(
        n11497) );
  OAI22_X2 U12234 ( .A1(n12278), .A2(n12776), .B1(n11498), .B2(n9507), .ZN(
        n11499) );
  AOI221_X2 U12235 ( .B1(n9511), .B2(n11801), .C1(n12780), .C2(n11500), .A(
        n11499), .ZN(n11504) );
  INV_X4 U12236 ( .A(n11501), .ZN(n12642) );
  NAND2_X2 U12237 ( .A1(n12642), .A2(n9508), .ZN(n11503) );
  OAI22_X2 U12238 ( .A1(n11504), .A2(n12772), .B1(n6806), .B2(n12058), .ZN(
        n11505) );
  INV_X4 U12239 ( .A(n11507), .ZN(n12268) );
  NOR2_X2 U12240 ( .A1(n11757), .A2(n12776), .ZN(n11508) );
  NOR2_X2 U12241 ( .A1(n12780), .A2(n11508), .ZN(n11509) );
  MUX2_X2 U12242 ( .A(n12793), .B(n9479), .S(n11510), .Z(n11511) );
  NOR2_X2 U12243 ( .A1(n9513), .A2(n11511), .ZN(n11512) );
  OAI22_X2 U12244 ( .A1(n12785), .A2(n12085), .B1(n11513), .B2(n11512), .ZN(
        n11514) );
  AOI221_X2 U12245 ( .B1(pipeline_alu_N69), .B2(n6813), .C1(pipeline_alu_N263), 
        .C2(n6812), .A(n11514), .ZN(n11515) );
  NAND2_X2 U12246 ( .A1(n11516), .A2(n11515), .ZN(dmem_haddr[10]) );
  MUX2_X2 U12247 ( .A(pipeline_alu_out_WB[10]), .B(dmem_haddr[10]), .S(n9524), 
        .Z(n5834) );
  OAI22_X2 U12248 ( .A1(n12805), .A2(n11517), .B1(n545), .B2(n9498), .ZN(
        n11518) );
  AOI221_X2 U12249 ( .B1(n12668), .B2(n11519), .C1(pipeline_alu_out_WB[10]), 
        .C2(n12809), .A(n11518), .ZN(n11520) );
  INV_X4 U12250 ( .A(n11520), .ZN(n5802) );
  NAND2_X2 U12251 ( .A1(pipeline_csr_N311), .A2(n6750), .ZN(n11521) );
  OAI221_X2 U12252 ( .B1(n11527), .B2(n6705), .C1(n1493), .C2(n6687), .A(
        n11521), .ZN(n5865) );
  OAI22_X2 U12253 ( .A1(n6659), .A2(n11527), .B1(n1265), .B2(n6689), .ZN(n6091) );
  OAI22_X2 U12254 ( .A1(n6702), .A2(n11527), .B1(n10974), .B2(n9529), .ZN(
        n6166) );
  OAI22_X2 U12255 ( .A1(n6688), .A2(n11527), .B1(n1171), .B2(n3689), .ZN(n6134) );
  INV_X4 U12256 ( .A(pipeline_csr_N658), .ZN(n11522) );
  OAI22_X2 U12257 ( .A1(n12255), .A2(n11529), .B1(n6821), .B2(n11522), .ZN(
        pipeline_csr_N1898) );
  OAI22_X2 U12258 ( .A1(n6703), .A2(n11527), .B1(n10977), .B2(n3683), .ZN(
        n6071) );
  NAND2_X2 U12259 ( .A1(pipeline_csr_N818), .A2(n9476), .ZN(n11523) );
  OAI221_X2 U12260 ( .B1(n11527), .B2(n6704), .C1(n10978), .C2(n12352), .A(
        n11523), .ZN(n6004) );
  INV_X4 U12261 ( .A(pipeline_csr_N754), .ZN(n11524) );
  OAI22_X2 U12262 ( .A1(n9492), .A2(n11529), .B1(n9403), .B2(n11524), .ZN(
        pipeline_csr_N1994) );
  INV_X4 U12263 ( .A(pipeline_csr_N690), .ZN(n11525) );
  OAI22_X2 U12264 ( .A1(n9469), .A2(n11529), .B1(n9404), .B2(n11525), .ZN(
        pipeline_csr_N1930) );
  NAND2_X2 U12265 ( .A1(pipeline_csr_N786), .A2(n12346), .ZN(n11526) );
  OAI221_X2 U12266 ( .B1(n11527), .B2(n12347), .C1(n10980), .C2(n12349), .A(
        n11526), .ZN(n6036) );
  INV_X4 U12267 ( .A(pipeline_csr_N722), .ZN(n11528) );
  OAI22_X2 U12268 ( .A1(n12612), .A2(n11529), .B1(n9406), .B2(n11528), .ZN(
        pipeline_csr_N1962) );
  OAI22_X2 U12269 ( .A1(n7201), .A2(n6691), .B1(n428), .B2(n9523), .ZN(n6344)
         );
  INV_X4 U12270 ( .A(n11577), .ZN(n11835) );
  MUX2_X2 U12271 ( .A(n11834), .B(n11835), .S(n9399), .Z(n12169) );
  INV_X4 U12272 ( .A(n12169), .ZN(n11583) );
  INV_X4 U12273 ( .A(n11576), .ZN(n11836) );
  NAND2_X2 U12274 ( .A1(n11836), .A2(n9508), .ZN(n11530) );
  INV_X4 U12275 ( .A(n12127), .ZN(n11539) );
  INV_X4 U12276 ( .A(n11830), .ZN(n12164) );
  NAND2_X2 U12277 ( .A1(n9511), .A2(n11829), .ZN(n11531) );
  NOR2_X2 U12278 ( .A1(pipeline_alu_src_b[19]), .A2(n12357), .ZN(n11533) );
  NOR2_X2 U12279 ( .A1(n9513), .A2(n11533), .ZN(n11536) );
  OAI221_X2 U12280 ( .B1(n11548), .B2(n11536), .C1(n11535), .C2(n11534), .A(
        n12659), .ZN(n11537) );
  AOI221_X2 U12281 ( .B1(n11539), .B2(n12165), .C1(n12172), .C2(n11538), .A(
        n11537), .ZN(n11554) );
  NAND2_X2 U12282 ( .A1(n12780), .A2(n7006), .ZN(n11772) );
  INV_X4 U12283 ( .A(n11772), .ZN(n11541) );
  NOR2_X2 U12284 ( .A1(n11835), .A2(n12645), .ZN(n11540) );
  NOR2_X2 U12285 ( .A1(n11541), .A2(n11540), .ZN(n11542) );
  OAI221_X2 U12286 ( .B1(n11836), .B2(n9507), .C1(n11543), .C2(n9509), .A(
        n11542), .ZN(n11544) );
  INV_X4 U12287 ( .A(n11544), .ZN(n12128) );
  AOI221_X2 U12288 ( .B1(n9471), .B2(n11547), .C1(n12276), .C2(n11546), .A(
        n11545), .ZN(n12161) );
  INV_X4 U12289 ( .A(n12161), .ZN(n12581) );
  MUX2_X2 U12290 ( .A(n12355), .B(n12357), .S(n11548), .Z(n11549) );
  NAND2_X2 U12291 ( .A1(n11549), .A2(n9512), .ZN(n11550) );
  NAND2_X2 U12292 ( .A1(n11550), .A2(pipeline_alu_src_b[19]), .ZN(n11551) );
  OAI221_X2 U12293 ( .B1(n12128), .B2(n12639), .C1(n12581), .C2(n12182), .A(
        n11551), .ZN(n11552) );
  AOI221_X2 U12294 ( .B1(pipeline_alu_N78), .B2(n6813), .C1(pipeline_alu_N272), 
        .C2(n6812), .A(n11552), .ZN(n11553) );
  NAND2_X2 U12295 ( .A1(n11554), .A2(n11553), .ZN(dmem_haddr[19]) );
  MUX2_X2 U12296 ( .A(pipeline_alu_out_WB[19]), .B(dmem_haddr[19]), .S(n9522), 
        .Z(n5825) );
  OAI22_X2 U12297 ( .A1(n12805), .A2(n11555), .B1(n554), .B2(n9498), .ZN(
        n11556) );
  AOI221_X2 U12298 ( .B1(n12668), .B2(n11557), .C1(pipeline_alu_out_WB[19]), 
        .C2(n12809), .A(n11556), .ZN(n11558) );
  INV_X4 U12299 ( .A(n11558), .ZN(n5793) );
  NAND2_X2 U12300 ( .A1(pipeline_csr_N320), .A2(n6750), .ZN(n11559) );
  OAI221_X2 U12301 ( .B1(n11565), .B2(n6705), .C1(n1502), .C2(n6687), .A(
        n11559), .ZN(n5856) );
  OAI22_X2 U12302 ( .A1(n6659), .A2(n11565), .B1(n1274), .B2(n6689), .ZN(n6100) );
  OAI22_X2 U12303 ( .A1(n6702), .A2(n11565), .B1(n10947), .B2(n9529), .ZN(
        n6157) );
  OAI22_X2 U12304 ( .A1(n6688), .A2(n11565), .B1(n1180), .B2(n3689), .ZN(n6125) );
  INV_X4 U12305 ( .A(pipeline_csr_N667), .ZN(n11560) );
  OAI22_X2 U12306 ( .A1(n12255), .A2(n11567), .B1(n6821), .B2(n11560), .ZN(
        pipeline_csr_N1907) );
  OAI22_X2 U12307 ( .A1(n6703), .A2(n11565), .B1(n10950), .B2(n3683), .ZN(
        n6062) );
  NAND2_X2 U12308 ( .A1(pipeline_csr_N827), .A2(n9476), .ZN(n11561) );
  OAI221_X2 U12309 ( .B1(n11565), .B2(n6704), .C1(n10951), .C2(n12352), .A(
        n11561), .ZN(n5995) );
  INV_X4 U12310 ( .A(pipeline_csr_N763), .ZN(n11562) );
  OAI22_X2 U12311 ( .A1(n9492), .A2(n11567), .B1(n9403), .B2(n11562), .ZN(
        pipeline_csr_N2003) );
  INV_X4 U12312 ( .A(pipeline_csr_N699), .ZN(n11563) );
  OAI22_X2 U12313 ( .A1(n9469), .A2(n11567), .B1(n9404), .B2(n11563), .ZN(
        pipeline_csr_N1939) );
  NAND2_X2 U12314 ( .A1(pipeline_csr_N795), .A2(n12346), .ZN(n11564) );
  OAI221_X2 U12315 ( .B1(n11565), .B2(n12347), .C1(n10953), .C2(n12349), .A(
        n11564), .ZN(n6027) );
  INV_X4 U12316 ( .A(pipeline_csr_N731), .ZN(n11566) );
  OAI22_X2 U12317 ( .A1(n12612), .A2(n11567), .B1(n9405), .B2(n11566), .ZN(
        pipeline_csr_N1971) );
  OAI22_X2 U12318 ( .A1(n7194), .A2(n6691), .B1(n446), .B2(n9523), .ZN(n6353)
         );
  NAND2_X2 U12319 ( .A1(n9479), .A2(n11589), .ZN(n11568) );
  NAND2_X2 U12320 ( .A1(n11568), .A2(n9512), .ZN(n11582) );
  INV_X4 U12321 ( .A(n12135), .ZN(n11874) );
  OAI22_X2 U12322 ( .A1(n11874), .A2(n12776), .B1(n12133), .B2(n9507), .ZN(
        n11575) );
  AOI221_X2 U12323 ( .B1(n9511), .B2(n11876), .C1(n12780), .C2(n11576), .A(
        n11575), .ZN(n11580) );
  NAND2_X2 U12324 ( .A1(n9510), .A2(n11577), .ZN(n11578) );
  OAI22_X2 U12325 ( .A1(n11580), .A2(n12772), .B1(n6746), .B2(n11579), .ZN(
        n11581) );
  NOR2_X2 U12326 ( .A1(n12776), .A2(n11829), .ZN(n11585) );
  NOR2_X2 U12327 ( .A1(n12780), .A2(n11585), .ZN(n11586) );
  MUX2_X2 U12328 ( .A(n12793), .B(n9479), .S(n6613), .Z(n11587) );
  NOR2_X2 U12329 ( .A1(n9513), .A2(n11587), .ZN(n11588) );
  OAI22_X2 U12330 ( .A1(n12785), .A2(n12160), .B1(n11589), .B2(n11588), .ZN(
        n11590) );
  AOI221_X2 U12331 ( .B1(pipeline_alu_N70), .B2(n6813), .C1(pipeline_alu_N264), 
        .C2(n6812), .A(n11590), .ZN(n11591) );
  NAND2_X2 U12332 ( .A1(n11592), .A2(n11591), .ZN(dmem_haddr[11]) );
  MUX2_X2 U12333 ( .A(pipeline_alu_out_WB[11]), .B(dmem_haddr[11]), .S(n9523), 
        .Z(n5833) );
  OAI22_X2 U12334 ( .A1(n12805), .A2(n11593), .B1(n546), .B2(n9498), .ZN(
        n11594) );
  AOI221_X2 U12335 ( .B1(n12668), .B2(n11595), .C1(pipeline_alu_out_WB[11]), 
        .C2(n12809), .A(n11594), .ZN(n11596) );
  INV_X4 U12336 ( .A(n11596), .ZN(n5801) );
  NAND2_X2 U12337 ( .A1(pipeline_csr_N312), .A2(n6750), .ZN(n11597) );
  OAI221_X2 U12338 ( .B1(n11603), .B2(n6705), .C1(n1494), .C2(n6687), .A(
        n11597), .ZN(n5864) );
  OAI22_X2 U12339 ( .A1(n6659), .A2(n11603), .B1(n1266), .B2(n6689), .ZN(n6092) );
  OAI22_X2 U12340 ( .A1(n6702), .A2(n11603), .B1(n10920), .B2(n9529), .ZN(
        n6165) );
  OAI22_X2 U12341 ( .A1(n6688), .A2(n11603), .B1(n1172), .B2(n3689), .ZN(n6133) );
  INV_X4 U12342 ( .A(pipeline_csr_N659), .ZN(n11598) );
  OAI22_X2 U12343 ( .A1(n12255), .A2(n11605), .B1(n6821), .B2(n11598), .ZN(
        pipeline_csr_N1899) );
  OAI22_X2 U12344 ( .A1(n6703), .A2(n11603), .B1(n10923), .B2(n3683), .ZN(
        n6070) );
  NAND2_X2 U12345 ( .A1(pipeline_csr_N819), .A2(n12350), .ZN(n11599) );
  OAI221_X2 U12346 ( .B1(n11603), .B2(n6704), .C1(n10924), .C2(n12352), .A(
        n11599), .ZN(n6003) );
  INV_X4 U12347 ( .A(pipeline_csr_N755), .ZN(n11600) );
  OAI22_X2 U12348 ( .A1(n9492), .A2(n11605), .B1(n9403), .B2(n11600), .ZN(
        pipeline_csr_N1995) );
  INV_X4 U12349 ( .A(pipeline_csr_N691), .ZN(n11601) );
  OAI22_X2 U12350 ( .A1(n9469), .A2(n11605), .B1(n12257), .B2(n11601), .ZN(
        pipeline_csr_N1931) );
  NAND2_X2 U12351 ( .A1(pipeline_csr_N787), .A2(n12346), .ZN(n11602) );
  OAI221_X2 U12352 ( .B1(n11603), .B2(n12347), .C1(n10926), .C2(n12349), .A(
        n11602), .ZN(n6035) );
  INV_X4 U12353 ( .A(pipeline_csr_N723), .ZN(n11604) );
  OAI22_X2 U12354 ( .A1(n12612), .A2(n11605), .B1(n9405), .B2(n11604), .ZN(
        pipeline_csr_N1963) );
  OAI22_X2 U12355 ( .A1(n7200), .A2(n6691), .B1(n430), .B2(n9524), .ZN(n6345)
         );
  INV_X4 U12356 ( .A(n11952), .ZN(n11608) );
  NAND2_X2 U12357 ( .A1(n9511), .A2(n12208), .ZN(n11606) );
  OAI221_X2 U12358 ( .B1(n11608), .B2(n9507), .C1(n11607), .C2(n9509), .A(
        n11606), .ZN(n11616) );
  INV_X4 U12359 ( .A(n11946), .ZN(n11650) );
  NAND2_X2 U12360 ( .A1(n11653), .A2(n9511), .ZN(n11609) );
  MUX2_X2 U12361 ( .A(n11610), .B(n11944), .S(n9399), .Z(n12786) );
  NOR2_X2 U12362 ( .A1(n9513), .A2(n11611), .ZN(n11612) );
  OAI221_X2 U12363 ( .B1(n12786), .B2(n11613), .C1(n6925), .C2(n11612), .A(
        n12659), .ZN(n11614) );
  AOI221_X2 U12364 ( .B1(n12165), .B2(n11616), .C1(n12172), .C2(n11615), .A(
        n11614), .ZN(n11626) );
  INV_X4 U12365 ( .A(n11616), .ZN(n12795) );
  NAND4_X2 U12366 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n12219) );
  INV_X4 U12367 ( .A(n12219), .ZN(n11949) );
  MUX2_X2 U12368 ( .A(n12355), .B(n12357), .S(n6925), .Z(n11621) );
  NAND2_X2 U12369 ( .A1(n11621), .A2(n9512), .ZN(n11622) );
  NAND2_X2 U12370 ( .A1(n11622), .A2(pipeline_alu_src_b[20]), .ZN(n11623) );
  OAI221_X2 U12371 ( .B1(n6803), .B2(n12639), .C1(n11949), .C2(n12182), .A(
        n11623), .ZN(n11624) );
  AOI221_X2 U12372 ( .B1(pipeline_alu_N79), .B2(n6813), .C1(pipeline_alu_N273), 
        .C2(n6812), .A(n11624), .ZN(n11625) );
  NAND2_X2 U12373 ( .A1(n11626), .A2(n11625), .ZN(dmem_haddr[20]) );
  MUX2_X2 U12374 ( .A(pipeline_alu_out_WB[20]), .B(dmem_haddr[20]), .S(n9524), 
        .Z(n5824) );
  OAI22_X2 U12375 ( .A1(n12805), .A2(n11627), .B1(n555), .B2(n9498), .ZN(
        n11628) );
  AOI221_X2 U12376 ( .B1(n12668), .B2(n11629), .C1(pipeline_alu_out_WB[20]), 
        .C2(n12809), .A(n11628), .ZN(n11630) );
  INV_X4 U12377 ( .A(n11630), .ZN(n5792) );
  NAND2_X2 U12378 ( .A1(pipeline_csr_N321), .A2(n6750), .ZN(n11631) );
  OAI221_X2 U12379 ( .B1(n11637), .B2(n6705), .C1(n1503), .C2(n6687), .A(
        n11631), .ZN(n5855) );
  OAI22_X2 U12380 ( .A1(n6659), .A2(n11637), .B1(n1275), .B2(n6689), .ZN(n6101) );
  OAI22_X2 U12381 ( .A1(n6703), .A2(n11637), .B1(n1243), .B2(n3683), .ZN(n6061) );
  INV_X4 U12382 ( .A(pipeline_csr_N764), .ZN(n11632) );
  OAI22_X2 U12383 ( .A1(n9492), .A2(n11639), .B1(n9403), .B2(n11632), .ZN(
        pipeline_csr_N2004) );
  NAND2_X2 U12384 ( .A1(pipeline_csr_N828), .A2(n12350), .ZN(n11633) );
  OAI221_X2 U12385 ( .B1(n11637), .B2(n6704), .C1(n1435), .C2(n12352), .A(
        n11633), .ZN(n5994) );
  OAI22_X2 U12386 ( .A1(n6702), .A2(n11637), .B1(n10891), .B2(n9529), .ZN(
        n6156) );
  OAI22_X2 U12387 ( .A1(n6688), .A2(n11637), .B1(n1181), .B2(n3689), .ZN(n6124) );
  INV_X4 U12388 ( .A(pipeline_csr_N732), .ZN(n11634) );
  OAI22_X2 U12389 ( .A1(n12612), .A2(n11639), .B1(n9406), .B2(n11634), .ZN(
        pipeline_csr_N1972) );
  INV_X4 U12390 ( .A(pipeline_csr_N668), .ZN(n11635) );
  OAI22_X2 U12391 ( .A1(n12255), .A2(n11639), .B1(n6821), .B2(n11635), .ZN(
        pipeline_csr_N1908) );
  NAND2_X2 U12392 ( .A1(pipeline_csr_N796), .A2(n12346), .ZN(n11636) );
  OAI221_X2 U12393 ( .B1(n11637), .B2(n12347), .C1(n10893), .C2(n12349), .A(
        n11636), .ZN(n6026) );
  INV_X4 U12394 ( .A(pipeline_csr_N700), .ZN(n11638) );
  OAI22_X2 U12395 ( .A1(n9469), .A2(n11639), .B1(n9404), .B2(n11638), .ZN(
        pipeline_csr_N1940) );
  OAI22_X2 U12396 ( .A1(n7187), .A2(n6691), .B1(n448), .B2(n9525), .ZN(n6354)
         );
  NAND2_X2 U12397 ( .A1(n9479), .A2(n11656), .ZN(n11640) );
  NAND2_X2 U12398 ( .A1(n11640), .A2(n9512), .ZN(n11649) );
  NAND2_X2 U12399 ( .A1(n9510), .A2(n12208), .ZN(n11642) );
  NAND2_X2 U12400 ( .A1(n11642), .A2(n11641), .ZN(n12226) );
  OAI22_X2 U12401 ( .A1(n12773), .A2(n9509), .B1(n11643), .B2(n9507), .ZN(
        n11644) );
  AOI221_X2 U12402 ( .B1(n9511), .B2(n11985), .C1(n12780), .C2(n11952), .A(
        n11644), .ZN(n11647) );
  INV_X4 U12403 ( .A(n12208), .ZN(n11646) );
  OAI22_X2 U12404 ( .A1(n11647), .A2(n12772), .B1(n11646), .B2(n11645), .ZN(
        n11648) );
  INV_X4 U12405 ( .A(n12786), .ZN(n11652) );
  NAND2_X2 U12406 ( .A1(n9508), .A2(n11650), .ZN(n11651) );
  MUX2_X2 U12407 ( .A(n12793), .B(n9479), .S(n6924), .Z(n11654) );
  NOR2_X2 U12408 ( .A1(n9513), .A2(n11654), .ZN(n11655) );
  OAI22_X2 U12409 ( .A1(n12785), .A2(n12218), .B1(n11656), .B2(n11655), .ZN(
        n11657) );
  AOI221_X2 U12410 ( .B1(pipeline_alu_N71), .B2(n6813), .C1(pipeline_alu_N265), 
        .C2(n6812), .A(n11657), .ZN(n11658) );
  NAND2_X2 U12411 ( .A1(n11659), .A2(n11658), .ZN(dmem_haddr[12]) );
  MUX2_X2 U12412 ( .A(pipeline_alu_out_WB[12]), .B(dmem_haddr[12]), .S(n9522), 
        .Z(n5832) );
  OAI22_X2 U12413 ( .A1(n12805), .A2(n11660), .B1(n547), .B2(n9498), .ZN(
        n11661) );
  AOI221_X2 U12414 ( .B1(n12668), .B2(n11662), .C1(pipeline_alu_out_WB[12]), 
        .C2(n12809), .A(n11661), .ZN(n11663) );
  INV_X4 U12415 ( .A(n11663), .ZN(n5800) );
  NAND2_X2 U12416 ( .A1(pipeline_csr_N313), .A2(n6750), .ZN(n11664) );
  OAI221_X2 U12417 ( .B1(n11670), .B2(n6705), .C1(n1495), .C2(n6687), .A(
        n11664), .ZN(n5863) );
  OAI22_X2 U12418 ( .A1(n6659), .A2(n11670), .B1(n1267), .B2(n6689), .ZN(n6093) );
  OAI22_X2 U12419 ( .A1(n6702), .A2(n11670), .B1(n10866), .B2(n9529), .ZN(
        n6164) );
  OAI22_X2 U12420 ( .A1(n6688), .A2(n11670), .B1(n1173), .B2(n3689), .ZN(n6132) );
  INV_X4 U12421 ( .A(pipeline_csr_N660), .ZN(n11665) );
  OAI22_X2 U12422 ( .A1(n12255), .A2(n11672), .B1(n6821), .B2(n11665), .ZN(
        pipeline_csr_N1900) );
  OAI22_X2 U12423 ( .A1(n6703), .A2(n11670), .B1(n10869), .B2(n3683), .ZN(
        n6069) );
  NAND2_X2 U12424 ( .A1(pipeline_csr_N820), .A2(n12350), .ZN(n11666) );
  OAI221_X2 U12425 ( .B1(n11670), .B2(n6704), .C1(n10870), .C2(n12352), .A(
        n11666), .ZN(n6002) );
  INV_X4 U12426 ( .A(pipeline_csr_N756), .ZN(n11667) );
  OAI22_X2 U12427 ( .A1(n9492), .A2(n11672), .B1(n9403), .B2(n11667), .ZN(
        pipeline_csr_N1996) );
  INV_X4 U12428 ( .A(pipeline_csr_N692), .ZN(n11668) );
  OAI22_X2 U12429 ( .A1(n9469), .A2(n11672), .B1(n9404), .B2(n11668), .ZN(
        pipeline_csr_N1932) );
  NAND2_X2 U12430 ( .A1(pipeline_csr_N788), .A2(n12346), .ZN(n11669) );
  OAI221_X2 U12431 ( .B1(n11670), .B2(n12347), .C1(n10872), .C2(n12349), .A(
        n11669), .ZN(n6034) );
  INV_X4 U12432 ( .A(pipeline_csr_N724), .ZN(n11671) );
  OAI22_X2 U12433 ( .A1(n12612), .A2(n11672), .B1(n9406), .B2(n11671), .ZN(
        pipeline_csr_N1964) );
  OAI22_X2 U12434 ( .A1(n7199), .A2(n6691), .B1(n432), .B2(n9523), .ZN(n6346)
         );
  INV_X4 U12435 ( .A(n11673), .ZN(n12362) );
  MUX2_X2 U12436 ( .A(n12362), .B(n12013), .S(n9399), .Z(n11674) );
  INV_X4 U12437 ( .A(n11733), .ZN(n11685) );
  INV_X4 U12438 ( .A(n12010), .ZN(n11677) );
  NAND2_X2 U12439 ( .A1(n11675), .A2(n9511), .ZN(n11676) );
  NOR2_X2 U12440 ( .A1(n9513), .A2(n11678), .ZN(n11682) );
  INV_X4 U12441 ( .A(n11679), .ZN(n12305) );
  OAI22_X2 U12442 ( .A1(n11681), .A2(n9509), .B1(n11680), .B2(n12774), .ZN(
        n11686) );
  OAI221_X2 U12443 ( .B1(n11693), .B2(n11682), .C1(n11725), .C2(n12089), .A(
        n12659), .ZN(n11683) );
  AOI221_X2 U12444 ( .B1(n11685), .B2(n12174), .C1(n12172), .C2(n11684), .A(
        n11683), .ZN(n11700) );
  INV_X4 U12445 ( .A(n11686), .ZN(n11688) );
  NAND2_X2 U12446 ( .A1(n9511), .A2(n12025), .ZN(n11687) );
  NAND3_X2 U12447 ( .A1(n11688), .A2(n11772), .A3(n11687), .ZN(n11728) );
  INV_X4 U12448 ( .A(n11728), .ZN(n11697) );
  NAND4_X2 U12449 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n12315) );
  INV_X4 U12450 ( .A(n12315), .ZN(n12016) );
  MUX2_X2 U12451 ( .A(n12355), .B(n12357), .S(n11693), .Z(n11694) );
  NAND2_X2 U12452 ( .A1(n11694), .A2(n9512), .ZN(n11695) );
  OAI221_X2 U12453 ( .B1(n11697), .B2(n12639), .C1(n12016), .C2(n12182), .A(
        n11696), .ZN(n11698) );
  AOI221_X2 U12454 ( .B1(pipeline_alu_N80), .B2(n6813), .C1(pipeline_alu_N274), 
        .C2(n6812), .A(n11698), .ZN(n11699) );
  NAND2_X2 U12455 ( .A1(n11700), .A2(n11699), .ZN(dmem_haddr[21]) );
  MUX2_X2 U12456 ( .A(pipeline_alu_out_WB[21]), .B(dmem_haddr[21]), .S(n9522), 
        .Z(n5823) );
  OAI22_X2 U12457 ( .A1(n12805), .A2(n11701), .B1(n556), .B2(n9498), .ZN(
        n11702) );
  AOI221_X2 U12458 ( .B1(n12668), .B2(n11703), .C1(pipeline_alu_out_WB[21]), 
        .C2(n12809), .A(n11702), .ZN(n11704) );
  INV_X4 U12459 ( .A(n11704), .ZN(n5791) );
  NAND2_X2 U12460 ( .A1(pipeline_csr_N322), .A2(n6750), .ZN(n11705) );
  OAI221_X2 U12461 ( .B1(n11711), .B2(n6705), .C1(n1504), .C2(n6687), .A(
        n11705), .ZN(n5854) );
  OAI22_X2 U12462 ( .A1(n6659), .A2(n11711), .B1(n1276), .B2(n6689), .ZN(n6102) );
  OAI22_X2 U12463 ( .A1(n6702), .A2(n11711), .B1(n10839), .B2(n9529), .ZN(
        n6155) );
  OAI22_X2 U12464 ( .A1(n6688), .A2(n11711), .B1(n1182), .B2(n3689), .ZN(n6123) );
  INV_X4 U12465 ( .A(pipeline_csr_N669), .ZN(n11706) );
  OAI22_X2 U12466 ( .A1(n12255), .A2(n11713), .B1(n6821), .B2(n11706), .ZN(
        pipeline_csr_N1909) );
  OAI22_X2 U12467 ( .A1(n6703), .A2(n11711), .B1(n10842), .B2(n3683), .ZN(
        n6060) );
  NAND2_X2 U12468 ( .A1(pipeline_csr_N829), .A2(n12350), .ZN(n11707) );
  OAI221_X2 U12469 ( .B1(n11711), .B2(n6704), .C1(n10843), .C2(n12352), .A(
        n11707), .ZN(n5993) );
  INV_X4 U12470 ( .A(pipeline_csr_N765), .ZN(n11708) );
  OAI22_X2 U12471 ( .A1(n9492), .A2(n11713), .B1(n9403), .B2(n11708), .ZN(
        pipeline_csr_N2005) );
  INV_X4 U12472 ( .A(pipeline_csr_N701), .ZN(n11709) );
  OAI22_X2 U12473 ( .A1(n9469), .A2(n11713), .B1(n12257), .B2(n11709), .ZN(
        pipeline_csr_N1941) );
  NAND2_X2 U12474 ( .A1(pipeline_csr_N797), .A2(n12346), .ZN(n11710) );
  OAI221_X2 U12475 ( .B1(n11711), .B2(n12347), .C1(n10845), .C2(n12349), .A(
        n11710), .ZN(n6025) );
  INV_X4 U12476 ( .A(pipeline_csr_N733), .ZN(n11712) );
  OAI22_X2 U12477 ( .A1(n12612), .A2(n11713), .B1(n9405), .B2(n11712), .ZN(
        pipeline_csr_N1973) );
  OAI22_X2 U12478 ( .A1(n7203), .A2(n6691), .B1(n450), .B2(n9525), .ZN(n6355)
         );
  NAND2_X2 U12479 ( .A1(n9479), .A2(n11732), .ZN(n11714) );
  NAND2_X2 U12480 ( .A1(n11714), .A2(n9512), .ZN(n11729) );
  INV_X4 U12481 ( .A(n12371), .ZN(n11724) );
  NAND4_X2 U12482 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n12373) );
  INV_X4 U12483 ( .A(n12373), .ZN(n12054) );
  OAI22_X2 U12484 ( .A1(n6801), .A2(n12776), .B1(n12054), .B2(n9507), .ZN(
        n11723) );
  AOI221_X2 U12485 ( .B1(n9511), .B2(n11724), .C1(n12780), .C2(n12057), .A(
        n11723), .ZN(n11726) );
  OAI22_X2 U12486 ( .A1(n11726), .A2(n12772), .B1(n11725), .B2(n12058), .ZN(
        n11727) );
  MUX2_X2 U12487 ( .A(n12793), .B(n9479), .S(n6619), .Z(n11730) );
  NOR2_X2 U12488 ( .A1(n9513), .A2(n11730), .ZN(n11731) );
  OAI22_X2 U12489 ( .A1(n12785), .A2(n11733), .B1(n11732), .B2(n11731), .ZN(
        n11734) );
  AOI221_X2 U12490 ( .B1(pipeline_alu_N64), .B2(n6813), .C1(pipeline_alu_N258), 
        .C2(n6812), .A(n11734), .ZN(n11735) );
  NAND2_X2 U12491 ( .A1(n11736), .A2(n11735), .ZN(dmem_haddr[5]) );
  MUX2_X2 U12492 ( .A(pipeline_alu_out_WB[5]), .B(dmem_haddr[5]), .S(n9524), 
        .Z(n5839) );
  OAI22_X2 U12493 ( .A1(n12805), .A2(n11737), .B1(n540), .B2(n9498), .ZN(
        n11738) );
  AOI221_X2 U12494 ( .B1(n12668), .B2(n11739), .C1(pipeline_alu_out_WB[5]), 
        .C2(n12809), .A(n11738), .ZN(n11740) );
  INV_X4 U12495 ( .A(n11740), .ZN(n5807) );
  NAND3_X2 U12496 ( .A1(n12148), .A2(n13130), .A3(n11742), .ZN(n12159) );
  NAND2_X2 U12497 ( .A1(n12159), .A2(n13130), .ZN(n12817) );
  INV_X4 U12498 ( .A(n12817), .ZN(n11745) );
  INV_X4 U12499 ( .A(n11742), .ZN(n11743) );
  NAND2_X2 U12500 ( .A1(n11743), .A2(n13130), .ZN(n12820) );
  INV_X4 U12501 ( .A(n12396), .ZN(n11744) );
  NAND2_X2 U12502 ( .A1(n11744), .A2(n13130), .ZN(n12822) );
  NAND3_X2 U12503 ( .A1(n11745), .A2(n12820), .A3(n12822), .ZN(n12816) );
  INV_X4 U12504 ( .A(n12159), .ZN(n12811) );
  NAND2_X2 U12505 ( .A1(n12811), .A2(pipeline_ctrl_N82), .ZN(n11746) );
  OAI221_X2 U12506 ( .B1(n12821), .B2(n12816), .C1(n11752), .C2(n12820), .A(
        n11746), .ZN(n5980) );
  OAI22_X2 U12507 ( .A1(n11752), .A2(n6690), .B1(n1196), .B2(n6708), .ZN(n6203) );
  INV_X4 U12508 ( .A(pipeline_csr_N653), .ZN(n11747) );
  OAI22_X2 U12509 ( .A1(n12255), .A2(n11754), .B1(n6821), .B2(n11747), .ZN(
        pipeline_csr_N1893) );
  OAI22_X2 U12510 ( .A1(n6703), .A2(n11752), .B1(n1228), .B2(n3683), .ZN(n6076) );
  NAND2_X2 U12511 ( .A1(pipeline_csr_N813), .A2(n12350), .ZN(n11748) );
  OAI221_X2 U12512 ( .B1(n11752), .B2(n6704), .C1(n1420), .C2(n12352), .A(
        n11748), .ZN(n6009) );
  INV_X4 U12513 ( .A(pipeline_csr_N749), .ZN(n11749) );
  OAI22_X2 U12514 ( .A1(n12615), .A2(n11754), .B1(n9403), .B2(n11749), .ZN(
        pipeline_csr_N1989) );
  INV_X4 U12515 ( .A(pipeline_csr_N685), .ZN(n11750) );
  OAI22_X2 U12516 ( .A1(n9469), .A2(n11754), .B1(n9404), .B2(n11750), .ZN(
        pipeline_csr_N1925) );
  NAND2_X2 U12517 ( .A1(pipeline_csr_N781), .A2(n12346), .ZN(n11751) );
  OAI221_X2 U12518 ( .B1(n11752), .B2(n12347), .C1(n10785), .C2(n12349), .A(
        n11751), .ZN(n6041) );
  INV_X4 U12519 ( .A(pipeline_csr_N717), .ZN(n11753) );
  OAI22_X2 U12520 ( .A1(n12612), .A2(n11754), .B1(n9406), .B2(n11753), .ZN(
        pipeline_csr_N1957) );
  OAI22_X2 U12521 ( .A1(n6816), .A2(n6691), .B1(n418), .B2(n9524), .ZN(n6339)
         );
  MUX2_X2 U12522 ( .A(n12268), .B(n11755), .S(n9399), .Z(n11756) );
  INV_X4 U12523 ( .A(n11810), .ZN(n11768) );
  INV_X4 U12524 ( .A(n11757), .ZN(n11761) );
  NAND2_X2 U12525 ( .A1(n11758), .A2(n9511), .ZN(n11759) );
  NOR2_X2 U12526 ( .A1(n9513), .A2(n11762), .ZN(n11765) );
  OAI22_X2 U12527 ( .A1(n11764), .A2(n9509), .B1(n11763), .B2(n12774), .ZN(
        n11769) );
  OAI221_X2 U12528 ( .B1(n6624), .B2(n11765), .C1(n11802), .C2(n12089), .A(
        n12659), .ZN(n11766) );
  AOI221_X2 U12529 ( .B1(n11768), .B2(n12174), .C1(n12172), .C2(n11767), .A(
        n11766), .ZN(n11784) );
  INV_X4 U12530 ( .A(n11769), .ZN(n11773) );
  NAND2_X2 U12531 ( .A1(n9511), .A2(n11770), .ZN(n11771) );
  NAND3_X2 U12532 ( .A1(n11773), .A2(n11772), .A3(n11771), .ZN(n11805) );
  INV_X4 U12533 ( .A(n11805), .ZN(n11781) );
  MUX2_X2 U12534 ( .A(n12355), .B(n12357), .S(n6624), .Z(n11778) );
  NAND2_X2 U12535 ( .A1(n11778), .A2(n9512), .ZN(n11779) );
  NAND2_X2 U12536 ( .A1(n11779), .A2(pipeline_alu_src_b[22]), .ZN(n11780) );
  OAI221_X2 U12537 ( .B1(n11781), .B2(n12639), .C1(n6800), .C2(n12182), .A(
        n11780), .ZN(n11782) );
  AOI221_X2 U12538 ( .B1(pipeline_alu_N81), .B2(n6813), .C1(pipeline_alu_N275), 
        .C2(n6812), .A(n11782), .ZN(n11783) );
  NAND2_X2 U12539 ( .A1(n11784), .A2(n11783), .ZN(dmem_haddr[22]) );
  MUX2_X2 U12540 ( .A(pipeline_alu_out_WB[22]), .B(dmem_haddr[22]), .S(n9524), 
        .Z(n5822) );
  OAI22_X2 U12541 ( .A1(n12805), .A2(n11785), .B1(n557), .B2(n9498), .ZN(
        n11786) );
  AOI221_X2 U12542 ( .B1(n12668), .B2(n11787), .C1(pipeline_alu_out_WB[22]), 
        .C2(n12809), .A(n11786), .ZN(n11788) );
  INV_X4 U12543 ( .A(n11788), .ZN(n5790) );
  NAND2_X2 U12544 ( .A1(pipeline_csr_N323), .A2(n6750), .ZN(n11789) );
  OAI221_X2 U12545 ( .B1(n11795), .B2(n6705), .C1(n1505), .C2(n6687), .A(
        n11789), .ZN(n5853) );
  OAI22_X2 U12546 ( .A1(n6659), .A2(n11795), .B1(n1277), .B2(n6689), .ZN(n6103) );
  OAI22_X2 U12547 ( .A1(n6702), .A2(n11795), .B1(n10754), .B2(n9529), .ZN(
        n6154) );
  OAI22_X2 U12548 ( .A1(n6688), .A2(n11795), .B1(n1183), .B2(n3689), .ZN(n6122) );
  INV_X4 U12549 ( .A(pipeline_csr_N670), .ZN(n11790) );
  OAI22_X2 U12550 ( .A1(n12255), .A2(n11797), .B1(n6821), .B2(n11790), .ZN(
        pipeline_csr_N1910) );
  OAI22_X2 U12551 ( .A1(n6703), .A2(n11795), .B1(n10757), .B2(n3683), .ZN(
        n6059) );
  NAND2_X2 U12552 ( .A1(pipeline_csr_N830), .A2(n12350), .ZN(n11791) );
  OAI221_X2 U12553 ( .B1(n11795), .B2(n6704), .C1(n10758), .C2(n12352), .A(
        n11791), .ZN(n5992) );
  INV_X4 U12554 ( .A(pipeline_csr_N766), .ZN(n11792) );
  OAI22_X2 U12555 ( .A1(n12615), .A2(n11797), .B1(n9403), .B2(n11792), .ZN(
        pipeline_csr_N2006) );
  INV_X4 U12556 ( .A(pipeline_csr_N702), .ZN(n11793) );
  OAI22_X2 U12557 ( .A1(n9469), .A2(n11797), .B1(n12257), .B2(n11793), .ZN(
        pipeline_csr_N1942) );
  NAND2_X2 U12558 ( .A1(pipeline_csr_N798), .A2(n12346), .ZN(n11794) );
  OAI221_X2 U12559 ( .B1(n11795), .B2(n12347), .C1(n10760), .C2(n12349), .A(
        n11794), .ZN(n6024) );
  INV_X4 U12560 ( .A(pipeline_csr_N734), .ZN(n11796) );
  OAI22_X2 U12561 ( .A1(n12612), .A2(n11797), .B1(n9405), .B2(n11796), .ZN(
        pipeline_csr_N1974) );
  OAI22_X2 U12562 ( .A1(n7204), .A2(n6691), .B1(n452), .B2(n9525), .ZN(n6356)
         );
  NAND2_X2 U12563 ( .A1(n9479), .A2(n11809), .ZN(n11798) );
  NAND2_X2 U12564 ( .A1(n11798), .A2(n9512), .ZN(n11806) );
  OAI22_X2 U12565 ( .A1(n12272), .A2(n9509), .B1(n12278), .B2(n12774), .ZN(
        n11800) );
  AOI221_X2 U12566 ( .B1(n9511), .B2(n12281), .C1(n12780), .C2(n11801), .A(
        n11800), .ZN(n11803) );
  OAI22_X2 U12567 ( .A1(n11803), .A2(n12772), .B1(n11802), .B2(n12058), .ZN(
        n11804) );
  MUX2_X2 U12568 ( .A(n12793), .B(n9479), .S(n6604), .Z(n11807) );
  NOR2_X2 U12569 ( .A1(n9513), .A2(n11807), .ZN(n11808) );
  OAI22_X2 U12570 ( .A1(n12785), .A2(n11810), .B1(n11809), .B2(n11808), .ZN(
        n11811) );
  AOI221_X2 U12571 ( .B1(pipeline_alu_N65), .B2(n6813), .C1(pipeline_alu_N259), 
        .C2(n6812), .A(n11811), .ZN(n11812) );
  NAND2_X2 U12572 ( .A1(n11813), .A2(n11812), .ZN(dmem_haddr[6]) );
  MUX2_X2 U12573 ( .A(pipeline_alu_out_WB[6]), .B(dmem_haddr[6]), .S(n9522), 
        .Z(n5838) );
  OAI22_X2 U12574 ( .A1(n12805), .A2(n11814), .B1(n541), .B2(n9498), .ZN(
        n11815) );
  AOI221_X2 U12575 ( .B1(n12668), .B2(n11816), .C1(pipeline_alu_out_WB[6]), 
        .C2(n12809), .A(n11815), .ZN(n11817) );
  INV_X4 U12576 ( .A(n11817), .ZN(n5806) );
  NAND2_X2 U12577 ( .A1(pipeline_csr_N307), .A2(n6750), .ZN(n11818) );
  OAI221_X2 U12578 ( .B1(n11824), .B2(n6705), .C1(n1489), .C2(n6687), .A(
        n11818), .ZN(n5869) );
  OAI22_X2 U12579 ( .A1(n6659), .A2(n11824), .B1(n1261), .B2(n6689), .ZN(n6087) );
  OAI22_X2 U12580 ( .A1(n6703), .A2(n11824), .B1(n1229), .B2(n3683), .ZN(n6075) );
  INV_X4 U12581 ( .A(pipeline_csr_N686), .ZN(n11819) );
  OAI22_X2 U12582 ( .A1(n9469), .A2(n11826), .B1(n12257), .B2(n11819), .ZN(
        pipeline_csr_N1926) );
  NAND2_X2 U12583 ( .A1(pipeline_csr_N782), .A2(n9472), .ZN(n11820) );
  OAI221_X2 U12584 ( .B1(n11824), .B2(n12347), .C1(n1389), .C2(n12349), .A(
        n11820), .ZN(n6040) );
  OAI22_X2 U12585 ( .A1(n6702), .A2(n11824), .B1(n10731), .B2(n9529), .ZN(
        n6170) );
  OAI22_X2 U12586 ( .A1(n6688), .A2(n11824), .B1(n1167), .B2(n3689), .ZN(n6138) );
  INV_X4 U12587 ( .A(pipeline_csr_N718), .ZN(n11821) );
  OAI22_X2 U12588 ( .A1(n12612), .A2(n11826), .B1(n9405), .B2(n11821), .ZN(
        pipeline_csr_N1958) );
  INV_X4 U12589 ( .A(pipeline_csr_N654), .ZN(n11822) );
  OAI22_X2 U12590 ( .A1(n12255), .A2(n11826), .B1(n6821), .B2(n11822), .ZN(
        pipeline_csr_N1894) );
  NAND2_X2 U12591 ( .A1(pipeline_csr_N814), .A2(n12350), .ZN(n11823) );
  OAI221_X2 U12592 ( .B1(n11824), .B2(n6704), .C1(n10733), .C2(n12352), .A(
        n11823), .ZN(n6008) );
  INV_X4 U12593 ( .A(pipeline_csr_N750), .ZN(n11825) );
  OAI22_X2 U12594 ( .A1(n12615), .A2(n11826), .B1(n9403), .B2(n11825), .ZN(
        pipeline_csr_N1990) );
  OAI22_X2 U12595 ( .A1(n7186), .A2(n6691), .B1(n420), .B2(n9523), .ZN(n6340)
         );
  MUX2_X2 U12596 ( .A(n12126), .B(n11827), .S(n9399), .Z(n11828) );
  INV_X4 U12597 ( .A(n11886), .ZN(n11840) );
  INV_X4 U12598 ( .A(n11829), .ZN(n11832) );
  NAND2_X2 U12599 ( .A1(n11830), .A2(n9511), .ZN(n11831) );
  NOR2_X2 U12600 ( .A1(pipeline_alu_src_b[23]), .A2(n12357), .ZN(n11833) );
  NOR2_X2 U12601 ( .A1(n9513), .A2(n11833), .ZN(n11837) );
  INV_X4 U12602 ( .A(n11834), .ZN(n12576) );
  OAI22_X2 U12603 ( .A1(n11836), .A2(n9509), .B1(n11835), .B2(n12774), .ZN(
        n11841) );
  OAI221_X2 U12604 ( .B1(n11847), .B2(n11837), .C1(n11878), .C2(n12089), .A(
        n12659), .ZN(n11838) );
  AOI221_X2 U12605 ( .B1(n11840), .B2(n12174), .C1(n12172), .C2(n11839), .A(
        n11838), .ZN(n11854) );
  INV_X4 U12606 ( .A(n11841), .ZN(n11842) );
  NAND2_X2 U12607 ( .A1(n11842), .A2(n12027), .ZN(n11881) );
  INV_X4 U12608 ( .A(n11881), .ZN(n11851) );
  NAND4_X2 U12609 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n12579) );
  INV_X4 U12610 ( .A(n12579), .ZN(n12163) );
  MUX2_X2 U12611 ( .A(n12355), .B(n12357), .S(n11847), .Z(n11848) );
  NAND2_X2 U12612 ( .A1(n11848), .A2(n12783), .ZN(n11849) );
  NAND2_X2 U12613 ( .A1(n11849), .A2(pipeline_alu_src_b[23]), .ZN(n11850) );
  OAI221_X2 U12614 ( .B1(n11851), .B2(n12639), .C1(n12163), .C2(n12182), .A(
        n11850), .ZN(n11852) );
  AOI221_X2 U12615 ( .B1(pipeline_alu_N82), .B2(n6813), .C1(pipeline_alu_N276), 
        .C2(n6812), .A(n11852), .ZN(n11853) );
  NAND2_X2 U12616 ( .A1(n11854), .A2(n11853), .ZN(dmem_haddr[23]) );
  MUX2_X2 U12617 ( .A(pipeline_alu_out_WB[23]), .B(dmem_haddr[23]), .S(n9522), 
        .Z(n5821) );
  OAI22_X2 U12618 ( .A1(n12805), .A2(n11855), .B1(n558), .B2(n9498), .ZN(
        n11856) );
  AOI221_X2 U12619 ( .B1(n12668), .B2(n11857), .C1(pipeline_alu_out_WB[23]), 
        .C2(n12809), .A(n11856), .ZN(n11858) );
  INV_X4 U12620 ( .A(n11858), .ZN(n5789) );
  NAND2_X2 U12621 ( .A1(pipeline_csr_N324), .A2(n6750), .ZN(n11859) );
  OAI221_X2 U12622 ( .B1(n11867), .B2(n6705), .C1(n1506), .C2(n6687), .A(
        n11859), .ZN(n5852) );
  OAI22_X2 U12623 ( .A1(n6659), .A2(n11867), .B1(n1278), .B2(n6689), .ZN(n6104) );
  OAI22_X2 U12624 ( .A1(n6702), .A2(n11867), .B1(n10703), .B2(n9529), .ZN(
        n6153) );
  OAI22_X2 U12625 ( .A1(n6688), .A2(n11867), .B1(n1184), .B2(n9530), .ZN(n6121) );
  INV_X4 U12626 ( .A(pipeline_csr_N671), .ZN(n11860) );
  OAI22_X2 U12627 ( .A1(n12255), .A2(n11865), .B1(n6821), .B2(n11860), .ZN(
        pipeline_csr_N1911) );
  OAI22_X2 U12628 ( .A1(n6703), .A2(n11867), .B1(n10706), .B2(n3683), .ZN(
        n6058) );
  INV_X4 U12629 ( .A(pipeline_csr_N767), .ZN(n11861) );
  OAI22_X2 U12630 ( .A1(n12615), .A2(n11865), .B1(n9403), .B2(n11861), .ZN(
        pipeline_csr_N2007) );
  INV_X4 U12631 ( .A(pipeline_csr_N703), .ZN(n11862) );
  OAI22_X2 U12632 ( .A1(n9469), .A2(n11865), .B1(n9404), .B2(n11862), .ZN(
        pipeline_csr_N1943) );
  NAND2_X2 U12633 ( .A1(pipeline_csr_N831), .A2(n12350), .ZN(n11863) );
  OAI221_X2 U12634 ( .B1(n11867), .B2(n6704), .C1(n1438), .C2(n12352), .A(
        n11863), .ZN(n5991) );
  INV_X4 U12635 ( .A(pipeline_csr_N735), .ZN(n11864) );
  OAI22_X2 U12636 ( .A1(n12612), .A2(n11865), .B1(n9406), .B2(n11864), .ZN(
        pipeline_csr_N1975) );
  NAND2_X2 U12637 ( .A1(pipeline_csr_N799), .A2(n12346), .ZN(n11866) );
  OAI221_X2 U12638 ( .B1(n11867), .B2(n12347), .C1(n10708), .C2(n12349), .A(
        n11866), .ZN(n6023) );
  OAI22_X2 U12639 ( .A1(n7205), .A2(n6691), .B1(n454), .B2(n9524), .ZN(n6357)
         );
  NAND2_X2 U12640 ( .A1(n9479), .A2(n11885), .ZN(n11868) );
  NAND2_X2 U12641 ( .A1(n11868), .A2(n12783), .ZN(n11882) );
  OAI22_X2 U12642 ( .A1(n7082), .A2(n9509), .B1(n11874), .B2(n12774), .ZN(
        n11875) );
  AOI221_X2 U12643 ( .B1(n9511), .B2(n11877), .C1(n12780), .C2(n11876), .A(
        n11875), .ZN(n11879) );
  OAI22_X2 U12644 ( .A1(n11879), .A2(n12772), .B1(n11878), .B2(n12058), .ZN(
        n11880) );
  MUX2_X2 U12645 ( .A(n12793), .B(n9479), .S(n6610), .Z(n11883) );
  NOR2_X2 U12646 ( .A1(n9513), .A2(n11883), .ZN(n11884) );
  OAI22_X2 U12647 ( .A1(n12785), .A2(n11886), .B1(n11885), .B2(n11884), .ZN(
        n11887) );
  AOI221_X2 U12648 ( .B1(pipeline_alu_N66), .B2(n6813), .C1(pipeline_alu_N260), 
        .C2(n6812), .A(n11887), .ZN(n11888) );
  NAND2_X2 U12649 ( .A1(n11889), .A2(n11888), .ZN(dmem_haddr[7]) );
  MUX2_X2 U12650 ( .A(pipeline_alu_out_WB[7]), .B(dmem_haddr[7]), .S(n9522), 
        .Z(n5837) );
  OAI22_X2 U12651 ( .A1(n12805), .A2(n11890), .B1(n542), .B2(n9498), .ZN(
        n11891) );
  AOI221_X2 U12652 ( .B1(n12668), .B2(n11892), .C1(pipeline_alu_out_WB[7]), 
        .C2(n12809), .A(n11891), .ZN(n11893) );
  INV_X4 U12653 ( .A(n11893), .ZN(n5805) );
  NAND2_X2 U12654 ( .A1(pipeline_csr_N308), .A2(n6750), .ZN(n11894) );
  OAI221_X2 U12655 ( .B1(n1490), .B2(n6687), .C1(n11943), .C2(n6705), .A(
        n11894), .ZN(n5868) );
  OAI22_X2 U12656 ( .A1(n6702), .A2(n12198), .B1(n10465), .B2(n9529), .ZN(
        n6149) );
  OAI22_X2 U12657 ( .A1(n6702), .A2(n12120), .B1(n10541), .B2(n9529), .ZN(
        n6150) );
  OAI22_X2 U12658 ( .A1(n6702), .A2(n12052), .B1(n10595), .B2(n9529), .ZN(
        n6151) );
  OAI22_X2 U12659 ( .A1(n6702), .A2(n11982), .B1(n10649), .B2(n9529), .ZN(
        n6152) );
  OAI22_X2 U12660 ( .A1(n6702), .A2(n12082), .B1(n10568), .B2(n9529), .ZN(
        n6167) );
  OAI22_X2 U12661 ( .A1(n6702), .A2(n12007), .B1(n10620), .B2(n9529), .ZN(
        n6168) );
  OAI22_X2 U12662 ( .A1(n6702), .A2(n11943), .B1(n10677), .B2(n9529), .ZN(
        n6169) );
  NOR2_X2 U12663 ( .A1(htif_reset), .A2(n11943), .ZN(n11895) );
  MUX2_X2 U12664 ( .A(n6706), .B(n11895), .S(n6826), .Z(n11935) );
  XOR2_X2 U12665 ( .A(n6815), .B(pipeline_csr_mtimecmp[1]), .Z(n11903) );
  XOR2_X2 U12666 ( .A(n6850), .B(pipeline_csr_mtimecmp[2]), .Z(n11902) );
  XOR2_X2 U12667 ( .A(n6823), .B(pipeline_csr_mtimecmp[0]), .Z(n11901) );
  XOR2_X2 U12668 ( .A(pipeline_csr_mtimecmp[4]), .B(pipeline_csr_mtime_full[4]), .Z(n11899) );
  XOR2_X2 U12669 ( .A(pipeline_csr_mtime_full[3]), .B(pipeline_csr_mtimecmp[3]), .Z(n11898) );
  XOR2_X2 U12670 ( .A(pipeline_csr_mtimecmp[6]), .B(pipeline_csr_mtime_full[6]), .Z(n11897) );
  XOR2_X2 U12671 ( .A(pipeline_csr_mtimecmp[5]), .B(pipeline_csr_mtime_full[5]), .Z(n11896) );
  NOR4_X2 U12672 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11900) );
  NAND4_X2 U12673 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n11932) );
  XOR2_X2 U12674 ( .A(n6825), .B(pipeline_csr_mtimecmp[8]), .Z(n11911) );
  XOR2_X2 U12675 ( .A(n6860), .B(pipeline_csr_mtimecmp[9]), .Z(n11910) );
  XOR2_X2 U12676 ( .A(n6861), .B(pipeline_csr_mtimecmp[7]), .Z(n11909) );
  XOR2_X2 U12677 ( .A(pipeline_csr_mtimecmp[11]), .B(
        pipeline_csr_mtime_full[11]), .Z(n11907) );
  XOR2_X2 U12678 ( .A(pipeline_csr_mtimecmp[10]), .B(
        pipeline_csr_mtime_full[10]), .Z(n11906) );
  XOR2_X2 U12679 ( .A(pipeline_csr_mtimecmp[13]), .B(
        pipeline_csr_mtime_full[13]), .Z(n11905) );
  XOR2_X2 U12680 ( .A(pipeline_csr_mtimecmp[12]), .B(
        pipeline_csr_mtime_full[12]), .Z(n11904) );
  NOR4_X2 U12681 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11908) );
  NAND4_X2 U12682 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11931) );
  XOR2_X2 U12683 ( .A(n6865), .B(pipeline_csr_mtimecmp[15]), .Z(n11919) );
  XOR2_X2 U12684 ( .A(n6857), .B(pipeline_csr_mtimecmp[16]), .Z(n11918) );
  XOR2_X2 U12685 ( .A(n6858), .B(pipeline_csr_mtimecmp[14]), .Z(n11917) );
  XOR2_X2 U12686 ( .A(pipeline_csr_mtimecmp[18]), .B(
        pipeline_csr_mtime_full[18]), .Z(n11915) );
  XOR2_X2 U12687 ( .A(pipeline_csr_mtimecmp[17]), .B(
        pipeline_csr_mtime_full[17]), .Z(n11914) );
  XOR2_X2 U12688 ( .A(pipeline_csr_mtimecmp[20]), .B(
        pipeline_csr_mtime_full[20]), .Z(n11913) );
  XOR2_X2 U12689 ( .A(pipeline_csr_mtimecmp[19]), .B(
        pipeline_csr_mtime_full[19]), .Z(n11912) );
  NOR4_X2 U12690 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11916) );
  NAND4_X2 U12691 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11930) );
  XOR2_X2 U12692 ( .A(n6862), .B(pipeline_csr_mtimecmp[27]), .Z(n11928) );
  XOR2_X2 U12693 ( .A(pipeline_csr_mtimecmp[26]), .B(
        pipeline_csr_mtime_full[26]), .Z(n11921) );
  XOR2_X2 U12694 ( .A(pipeline_csr_mtimecmp[25]), .B(
        pipeline_csr_mtime_full[25]), .Z(n11920) );
  NOR2_X2 U12695 ( .A1(n11921), .A2(n11920), .ZN(n11927) );
  XOR2_X2 U12696 ( .A(pipeline_csr_mtimecmp[22]), .B(
        pipeline_csr_mtime_full[22]), .Z(n11925) );
  XOR2_X2 U12697 ( .A(pipeline_csr_mtimecmp[21]), .B(
        pipeline_csr_mtime_full[21]), .Z(n11924) );
  XOR2_X2 U12698 ( .A(pipeline_csr_mtimecmp[24]), .B(
        pipeline_csr_mtime_full[24]), .Z(n11923) );
  XOR2_X2 U12699 ( .A(pipeline_csr_mtimecmp[23]), .B(
        pipeline_csr_mtime_full[23]), .Z(n11922) );
  NOR4_X2 U12700 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11926) );
  NAND4_X2 U12701 ( .A1(n4147), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11929) );
  NOR4_X2 U12702 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n11933) );
  NOR3_X2 U12703 ( .A1(n11933), .A2(n9529), .A3(n6826), .ZN(n11934) );
  MUX2_X2 U12704 ( .A(n11935), .B(pipeline_csr_mip_7_), .S(n11934), .Z(n6366)
         );
  OAI22_X2 U12705 ( .A1(n6659), .A2(n11943), .B1(n1262), .B2(n6689), .ZN(n6088) );
  OAI22_X2 U12706 ( .A1(n6688), .A2(n11943), .B1(n1168), .B2(n9530), .ZN(n6137) );
  INV_X4 U12707 ( .A(pipeline_csr_N655), .ZN(n11936) );
  OAI22_X2 U12708 ( .A1(n12255), .A2(n11941), .B1(n6821), .B2(n11936), .ZN(
        pipeline_csr_N1895) );
  OAI22_X2 U12709 ( .A1(n6703), .A2(n11943), .B1(n10680), .B2(n3683), .ZN(
        n6074) );
  INV_X4 U12710 ( .A(pipeline_csr_N687), .ZN(n11937) );
  OAI22_X2 U12711 ( .A1(n9469), .A2(n11941), .B1(n9404), .B2(n11937), .ZN(
        pipeline_csr_N1927) );
  INV_X4 U12712 ( .A(pipeline_csr_N751), .ZN(n11938) );
  OAI22_X2 U12713 ( .A1(n12615), .A2(n11941), .B1(n9403), .B2(n11938), .ZN(
        pipeline_csr_N1991) );
  NAND2_X2 U12714 ( .A1(pipeline_csr_N815), .A2(n12350), .ZN(n11939) );
  OAI221_X2 U12715 ( .B1(n11943), .B2(n6704), .C1(n1422), .C2(n12352), .A(
        n11939), .ZN(n6007) );
  INV_X4 U12716 ( .A(pipeline_csr_N719), .ZN(n11940) );
  OAI22_X2 U12717 ( .A1(n12612), .A2(n11941), .B1(n9406), .B2(n11940), .ZN(
        pipeline_csr_N1959) );
  NAND2_X2 U12718 ( .A1(pipeline_csr_N783), .A2(n12346), .ZN(n11942) );
  OAI221_X2 U12719 ( .B1(n11943), .B2(n12347), .C1(n10682), .C2(n12349), .A(
        n11942), .ZN(n6039) );
  OAI22_X2 U12720 ( .A1(n7185), .A2(n6691), .B1(n422), .B2(n9524), .ZN(n6341)
         );
  NAND2_X2 U12721 ( .A1(n9508), .A2(n11944), .ZN(n11945) );
  INV_X4 U12722 ( .A(n11993), .ZN(n11957) );
  NAND2_X2 U12723 ( .A1(n11947), .A2(n9511), .ZN(n11948) );
  NOR2_X2 U12724 ( .A1(pipeline_alu_src_b[24]), .A2(n12357), .ZN(n11951) );
  NOR2_X2 U12725 ( .A1(n9513), .A2(n11951), .ZN(n11954) );
  MUX2_X2 U12726 ( .A(n12208), .B(n11952), .S(n9399), .Z(n11953) );
  OAI221_X2 U12727 ( .B1(n11962), .B2(n11954), .C1(n12089), .C2(n11986), .A(
        n12659), .ZN(n11955) );
  AOI221_X2 U12728 ( .B1(n11957), .B2(n12174), .C1(n12172), .C2(n11956), .A(
        n11955), .ZN(n11969) );
  NAND2_X2 U12729 ( .A1(n11986), .A2(n12027), .ZN(n11989) );
  INV_X4 U12730 ( .A(n11989), .ZN(n11966) );
  MUX2_X2 U12731 ( .A(n12355), .B(n12357), .S(n11962), .Z(n11963) );
  NAND2_X2 U12732 ( .A1(n11963), .A2(n12783), .ZN(n11964) );
  NAND2_X2 U12733 ( .A1(n11964), .A2(pipeline_alu_src_b[24]), .ZN(n11965) );
  OAI221_X2 U12734 ( .B1(n11966), .B2(n12639), .C1(n6804), .C2(n12182), .A(
        n11965), .ZN(n11967) );
  AOI221_X2 U12735 ( .B1(pipeline_alu_N83), .B2(n6813), .C1(pipeline_alu_N277), 
        .C2(n6812), .A(n11967), .ZN(n11968) );
  NAND2_X2 U12736 ( .A1(n11969), .A2(n11968), .ZN(dmem_haddr[24]) );
  MUX2_X2 U12737 ( .A(pipeline_alu_out_WB[24]), .B(dmem_haddr[24]), .S(n9523), 
        .Z(n5820) );
  OAI22_X2 U12738 ( .A1(n12805), .A2(n11970), .B1(n559), .B2(n9498), .ZN(
        n11971) );
  AOI221_X2 U12739 ( .B1(n12668), .B2(n11972), .C1(pipeline_alu_out_WB[24]), 
        .C2(n12809), .A(n11971), .ZN(n11973) );
  INV_X4 U12740 ( .A(n11973), .ZN(n5788) );
  NAND2_X2 U12741 ( .A1(pipeline_csr_N325), .A2(n6750), .ZN(n11974) );
  OAI221_X2 U12742 ( .B1(n11982), .B2(n6705), .C1(n1507), .C2(n6687), .A(
        n11974), .ZN(n5851) );
  OAI22_X2 U12743 ( .A1(n6659), .A2(n11982), .B1(n1279), .B2(n6689), .ZN(n6105) );
  OAI22_X2 U12744 ( .A1(n6688), .A2(n11982), .B1(n1185), .B2(n9530), .ZN(n6120) );
  INV_X4 U12745 ( .A(pipeline_csr_N672), .ZN(n11975) );
  OAI22_X2 U12746 ( .A1(n12255), .A2(n11980), .B1(n6821), .B2(n11975), .ZN(
        pipeline_csr_N1912) );
  OAI22_X2 U12747 ( .A1(n6703), .A2(n11982), .B1(n10652), .B2(n3683), .ZN(
        n6057) );
  INV_X4 U12748 ( .A(pipeline_csr_N768), .ZN(n11976) );
  OAI22_X2 U12749 ( .A1(n12615), .A2(n11980), .B1(n9403), .B2(n11976), .ZN(
        pipeline_csr_N2008) );
  INV_X4 U12750 ( .A(pipeline_csr_N704), .ZN(n11977) );
  OAI22_X2 U12751 ( .A1(n9469), .A2(n11980), .B1(n12257), .B2(n11977), .ZN(
        pipeline_csr_N1944) );
  NAND2_X2 U12752 ( .A1(pipeline_csr_N832), .A2(n12350), .ZN(n11978) );
  OAI221_X2 U12753 ( .B1(n11982), .B2(n6704), .C1(n1439), .C2(n12352), .A(
        n11978), .ZN(n5990) );
  INV_X4 U12754 ( .A(pipeline_csr_N736), .ZN(n11979) );
  OAI22_X2 U12755 ( .A1(n12612), .A2(n11980), .B1(n9405), .B2(n11979), .ZN(
        pipeline_csr_N1976) );
  NAND2_X2 U12756 ( .A1(pipeline_csr_N800), .A2(n12346), .ZN(n11981) );
  OAI221_X2 U12757 ( .B1(n11982), .B2(n12347), .C1(n10654), .C2(n12349), .A(
        n11981), .ZN(n6022) );
  OAI22_X2 U12758 ( .A1(n7206), .A2(n6691), .B1(n456), .B2(n9525), .ZN(n6358)
         );
  NAND2_X2 U12759 ( .A1(n9479), .A2(n9387), .ZN(n11983) );
  NAND2_X2 U12760 ( .A1(n11983), .A2(n12783), .ZN(n11990) );
  OAI22_X2 U12761 ( .A1(n12775), .A2(n12776), .B1(n12773), .B2(n9507), .ZN(
        n11984) );
  AOI221_X2 U12762 ( .B1(n9511), .B2(n12779), .C1(n12780), .C2(n11985), .A(
        n11984), .ZN(n11987) );
  OAI22_X2 U12763 ( .A1(n11987), .A2(n12772), .B1(n12058), .B2(n11986), .ZN(
        n11988) );
  MUX2_X2 U12764 ( .A(n12793), .B(n9479), .S(n9334), .Z(n11991) );
  NOR2_X2 U12765 ( .A1(n9513), .A2(n11991), .ZN(n11992) );
  OAI22_X2 U12766 ( .A1(n12785), .A2(n11993), .B1(n9387), .B2(n11992), .ZN(
        n11994) );
  AOI221_X2 U12767 ( .B1(pipeline_alu_N67), .B2(n6813), .C1(pipeline_alu_N261), 
        .C2(n6812), .A(n11994), .ZN(n11995) );
  NAND2_X2 U12768 ( .A1(n11996), .A2(n11995), .ZN(dmem_haddr[8]) );
  MUX2_X2 U12769 ( .A(pipeline_alu_out_WB[8]), .B(dmem_haddr[8]), .S(n9522), 
        .Z(n5836) );
  OAI22_X2 U12770 ( .A1(n12805), .A2(n11997), .B1(n543), .B2(n9498), .ZN(
        n11998) );
  AOI221_X2 U12771 ( .B1(n12668), .B2(n11999), .C1(pipeline_alu_out_WB[8]), 
        .C2(n12809), .A(n11998), .ZN(n12000) );
  INV_X4 U12772 ( .A(n12000), .ZN(n5804) );
  NAND2_X2 U12773 ( .A1(pipeline_csr_N309), .A2(n6750), .ZN(n12001) );
  OAI221_X2 U12774 ( .B1(n12007), .B2(n6705), .C1(n1491), .C2(n6687), .A(
        n12001), .ZN(n5867) );
  OAI22_X2 U12775 ( .A1(n6659), .A2(n12007), .B1(n1263), .B2(n6689), .ZN(n6089) );
  OAI22_X2 U12776 ( .A1(n6703), .A2(n12007), .B1(n1231), .B2(n3683), .ZN(n6073) );
  INV_X4 U12777 ( .A(pipeline_csr_N752), .ZN(n12002) );
  OAI22_X2 U12778 ( .A1(n9492), .A2(n12009), .B1(n9403), .B2(n12002), .ZN(
        pipeline_csr_N1992) );
  NAND2_X2 U12779 ( .A1(pipeline_csr_N816), .A2(n9476), .ZN(n12003) );
  OAI221_X2 U12780 ( .B1(n12007), .B2(n6704), .C1(n1423), .C2(n12352), .A(
        n12003), .ZN(n6006) );
  OAI22_X2 U12781 ( .A1(n6688), .A2(n12007), .B1(n1169), .B2(n9530), .ZN(n6136) );
  INV_X4 U12782 ( .A(pipeline_csr_N720), .ZN(n12004) );
  OAI22_X2 U12783 ( .A1(n12612), .A2(n12009), .B1(n9406), .B2(n12004), .ZN(
        pipeline_csr_N1960) );
  INV_X4 U12784 ( .A(pipeline_csr_N656), .ZN(n12005) );
  OAI22_X2 U12785 ( .A1(n12255), .A2(n12009), .B1(n6821), .B2(n12005), .ZN(
        pipeline_csr_N1896) );
  NAND2_X2 U12786 ( .A1(pipeline_csr_N784), .A2(n12346), .ZN(n12006) );
  OAI221_X2 U12787 ( .B1(n12007), .B2(n12347), .C1(n10622), .C2(n12349), .A(
        n12006), .ZN(n6038) );
  INV_X4 U12788 ( .A(pipeline_csr_N688), .ZN(n12008) );
  OAI22_X2 U12789 ( .A1(n9469), .A2(n12009), .B1(n9404), .B2(n12008), .ZN(
        pipeline_csr_N1928) );
  OAI22_X2 U12790 ( .A1(n7213), .A2(n6691), .B1(n424), .B2(n9523), .ZN(n6342)
         );
  NOR2_X2 U12791 ( .A1(n9509), .A2(n12010), .ZN(n12011) );
  NOR2_X2 U12792 ( .A1(n12780), .A2(n12011), .ZN(n12012) );
  INV_X4 U12793 ( .A(n12068), .ZN(n12024) );
  NAND2_X2 U12794 ( .A1(n12014), .A2(n9511), .ZN(n12015) );
  NOR2_X2 U12795 ( .A1(pipeline_alu_src_b[25]), .A2(n12357), .ZN(n12018) );
  NOR2_X2 U12796 ( .A1(n9513), .A2(n12018), .ZN(n12021) );
  NAND2_X2 U12797 ( .A1(n12305), .A2(n9508), .ZN(n12020) );
  NAND2_X2 U12798 ( .A1(n9510), .A2(n12019), .ZN(n12026) );
  OAI221_X2 U12799 ( .B1(n6607), .B2(n12021), .C1(n6802), .C2(n12089), .A(
        n12659), .ZN(n12022) );
  AOI221_X2 U12800 ( .B1(n12024), .B2(n12174), .C1(n12172), .C2(n12023), .A(
        n12022), .ZN(n12039) );
  NAND2_X2 U12801 ( .A1(n9508), .A2(n12025), .ZN(n12028) );
  NAND3_X2 U12802 ( .A1(n12028), .A2(n12027), .A3(n12026), .ZN(n12061) );
  INV_X4 U12803 ( .A(n12061), .ZN(n12036) );
  MUX2_X2 U12804 ( .A(n12355), .B(n12357), .S(n6607), .Z(n12033) );
  NAND2_X2 U12805 ( .A1(n12033), .A2(n9512), .ZN(n12034) );
  NAND2_X2 U12806 ( .A1(n12034), .A2(pipeline_alu_src_b[25]), .ZN(n12035) );
  OAI221_X2 U12807 ( .B1(n12036), .B2(n12639), .C1(n6805), .C2(n12182), .A(
        n12035), .ZN(n12037) );
  AOI221_X2 U12808 ( .B1(pipeline_alu_N84), .B2(n6813), .C1(pipeline_alu_N278), 
        .C2(n6812), .A(n12037), .ZN(n12038) );
  NAND2_X2 U12809 ( .A1(n12039), .A2(n12038), .ZN(dmem_haddr[25]) );
  MUX2_X2 U12810 ( .A(pipeline_alu_out_WB[25]), .B(dmem_haddr[25]), .S(n9524), 
        .Z(n5819) );
  OAI22_X2 U12811 ( .A1(n12805), .A2(n12040), .B1(n560), .B2(n9498), .ZN(
        n12041) );
  AOI221_X2 U12812 ( .B1(n12668), .B2(n12042), .C1(pipeline_alu_out_WB[25]), 
        .C2(n12809), .A(n12041), .ZN(n12043) );
  INV_X4 U12813 ( .A(n12043), .ZN(n5787) );
  NAND2_X2 U12814 ( .A1(pipeline_csr_N326), .A2(n6750), .ZN(n12044) );
  OAI221_X2 U12815 ( .B1(n12052), .B2(n6705), .C1(n1508), .C2(n6687), .A(
        n12044), .ZN(n5850) );
  OAI22_X2 U12816 ( .A1(n6659), .A2(n12052), .B1(n1280), .B2(n6689), .ZN(n6106) );
  OAI22_X2 U12817 ( .A1(n6688), .A2(n12052), .B1(n1186), .B2(n9530), .ZN(n6119) );
  INV_X4 U12818 ( .A(pipeline_csr_N673), .ZN(n12045) );
  OAI22_X2 U12819 ( .A1(n12255), .A2(n12050), .B1(n6821), .B2(n12045), .ZN(
        pipeline_csr_N1913) );
  OAI22_X2 U12820 ( .A1(n6703), .A2(n12052), .B1(n10598), .B2(n3683), .ZN(
        n6056) );
  INV_X4 U12821 ( .A(pipeline_csr_N769), .ZN(n12046) );
  OAI22_X2 U12822 ( .A1(n12615), .A2(n12050), .B1(n9403), .B2(n12046), .ZN(
        pipeline_csr_N2009) );
  INV_X4 U12823 ( .A(pipeline_csr_N705), .ZN(n12047) );
  OAI22_X2 U12824 ( .A1(n9469), .A2(n12050), .B1(n12257), .B2(n12047), .ZN(
        pipeline_csr_N1945) );
  NAND2_X2 U12825 ( .A1(pipeline_csr_N833), .A2(n9476), .ZN(n12048) );
  OAI221_X2 U12826 ( .B1(n12052), .B2(n6704), .C1(n1440), .C2(n12352), .A(
        n12048), .ZN(n5989) );
  INV_X4 U12827 ( .A(pipeline_csr_N737), .ZN(n12049) );
  OAI22_X2 U12828 ( .A1(n12612), .A2(n12050), .B1(n9405), .B2(n12049), .ZN(
        pipeline_csr_N1977) );
  NAND2_X2 U12829 ( .A1(pipeline_csr_N801), .A2(n12346), .ZN(n12051) );
  OAI221_X2 U12830 ( .B1(n12052), .B2(n12347), .C1(n10600), .C2(n12349), .A(
        n12051), .ZN(n6021) );
  OAI22_X2 U12831 ( .A1(n7207), .A2(n6691), .B1(n458), .B2(n9524), .ZN(n6359)
         );
  NAND2_X2 U12832 ( .A1(n9479), .A2(n12067), .ZN(n12053) );
  NAND2_X2 U12833 ( .A1(n12053), .A2(n12783), .ZN(n12063) );
  OAI22_X2 U12834 ( .A1(n12054), .A2(n9509), .B1(n12371), .B2(n12774), .ZN(
        n12055) );
  AOI221_X2 U12835 ( .B1(n9511), .B2(n12057), .C1(n12780), .C2(n12056), .A(
        n12055), .ZN(n12059) );
  OAI22_X2 U12836 ( .A1(n12059), .A2(n12772), .B1(n6802), .B2(n12058), .ZN(
        n12060) );
  AOI221_X2 U12837 ( .B1(n12063), .B2(n6973), .C1(n12062), .C2(n12061), .A(
        n12060), .ZN(n12071) );
  MUX2_X2 U12838 ( .A(n12793), .B(n9479), .S(n12064), .Z(n12065) );
  NOR2_X2 U12839 ( .A1(n9513), .A2(n12065), .ZN(n12066) );
  OAI22_X2 U12840 ( .A1(n12785), .A2(n12068), .B1(n12067), .B2(n12066), .ZN(
        n12069) );
  AOI221_X2 U12841 ( .B1(pipeline_alu_N68), .B2(n6813), .C1(pipeline_alu_N262), 
        .C2(n6812), .A(n12069), .ZN(n12070) );
  NAND2_X2 U12842 ( .A1(n12071), .A2(n12070), .ZN(dmem_haddr[9]) );
  MUX2_X2 U12843 ( .A(pipeline_alu_out_WB[9]), .B(dmem_haddr[9]), .S(n9523), 
        .Z(n5835) );
  OAI22_X2 U12844 ( .A1(n12805), .A2(n12072), .B1(n544), .B2(n9498), .ZN(
        n12073) );
  AOI221_X2 U12845 ( .B1(n12668), .B2(n12074), .C1(pipeline_alu_out_WB[9]), 
        .C2(n12809), .A(n12073), .ZN(n12075) );
  INV_X4 U12846 ( .A(n12075), .ZN(n5803) );
  NAND2_X2 U12847 ( .A1(pipeline_csr_N310), .A2(n6750), .ZN(n12076) );
  OAI221_X2 U12848 ( .B1(n12082), .B2(n6705), .C1(n1492), .C2(n6687), .A(
        n12076), .ZN(n5866) );
  OAI22_X2 U12849 ( .A1(n6659), .A2(n12082), .B1(n1264), .B2(n6689), .ZN(n6090) );
  OAI22_X2 U12850 ( .A1(n6688), .A2(n12082), .B1(n1170), .B2(n3689), .ZN(n6135) );
  INV_X4 U12851 ( .A(pipeline_csr_N657), .ZN(n12077) );
  OAI22_X2 U12852 ( .A1(n12255), .A2(n12084), .B1(n6821), .B2(n12077), .ZN(
        pipeline_csr_N1897) );
  OAI22_X2 U12853 ( .A1(n6703), .A2(n12082), .B1(n10571), .B2(n3683), .ZN(
        n6072) );
  NAND2_X2 U12854 ( .A1(pipeline_csr_N817), .A2(n12350), .ZN(n12078) );
  OAI221_X2 U12855 ( .B1(n12082), .B2(n6704), .C1(n10572), .C2(n12352), .A(
        n12078), .ZN(n6005) );
  INV_X4 U12856 ( .A(pipeline_csr_N753), .ZN(n12079) );
  OAI22_X2 U12857 ( .A1(n12615), .A2(n12084), .B1(n9403), .B2(n12079), .ZN(
        pipeline_csr_N1993) );
  INV_X4 U12858 ( .A(pipeline_csr_N689), .ZN(n12080) );
  OAI22_X2 U12859 ( .A1(n9469), .A2(n12084), .B1(n12257), .B2(n12080), .ZN(
        pipeline_csr_N1929) );
  NAND2_X2 U12860 ( .A1(pipeline_csr_N785), .A2(n12346), .ZN(n12081) );
  OAI221_X2 U12861 ( .B1(n12082), .B2(n12347), .C1(n10574), .C2(n12349), .A(
        n12081), .ZN(n6037) );
  INV_X4 U12862 ( .A(pipeline_csr_N721), .ZN(n12083) );
  OAI22_X2 U12863 ( .A1(n12612), .A2(n12084), .B1(n9405), .B2(n12083), .ZN(
        pipeline_csr_N1961) );
  OAI22_X2 U12864 ( .A1(n7202), .A2(n6691), .B1(n426), .B2(n9525), .ZN(n6343)
         );
  INV_X4 U12865 ( .A(n12085), .ZN(n12093) );
  NAND2_X2 U12866 ( .A1(n12647), .A2(n9511), .ZN(n12086) );
  NOR2_X2 U12867 ( .A1(n9513), .A2(n12088), .ZN(n12090) );
  AOI221_X2 U12868 ( .B1(n12093), .B2(n12174), .C1(n12172), .C2(n12092), .A(
        n12091), .ZN(n12107) );
  INV_X4 U12869 ( .A(n12094), .ZN(n12104) );
  NAND4_X2 U12870 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12648) );
  INV_X4 U12871 ( .A(n12648), .ZN(n12103) );
  MUX2_X2 U12872 ( .A(n12355), .B(n12357), .S(n12099), .Z(n12100) );
  NAND2_X2 U12873 ( .A1(n12100), .A2(n12783), .ZN(n12101) );
  NAND2_X2 U12874 ( .A1(n12101), .A2(pipeline_alu_src_b[26]), .ZN(n12102) );
  OAI221_X2 U12875 ( .B1(n12104), .B2(n12639), .C1(n12103), .C2(n12182), .A(
        n12102), .ZN(n12105) );
  AOI221_X2 U12876 ( .B1(pipeline_alu_N85), .B2(n6813), .C1(pipeline_alu_N279), 
        .C2(n6812), .A(n12105), .ZN(n12106) );
  NAND2_X2 U12877 ( .A1(n12107), .A2(n12106), .ZN(dmem_haddr[26]) );
  MUX2_X2 U12878 ( .A(pipeline_alu_out_WB[26]), .B(dmem_haddr[26]), .S(n9525), 
        .Z(n5818) );
  OAI22_X2 U12879 ( .A1(n12805), .A2(n12108), .B1(n561), .B2(n9498), .ZN(
        n12109) );
  AOI221_X2 U12880 ( .B1(n12668), .B2(n12110), .C1(pipeline_alu_out_WB[26]), 
        .C2(n12809), .A(n12109), .ZN(n12111) );
  INV_X4 U12881 ( .A(n12111), .ZN(n5786) );
  NAND2_X2 U12882 ( .A1(pipeline_csr_N327), .A2(n6750), .ZN(n12112) );
  OAI221_X2 U12883 ( .B1(n12120), .B2(n6705), .C1(n1509), .C2(n6687), .A(
        n12112), .ZN(n5849) );
  OAI22_X2 U12884 ( .A1(n6659), .A2(n12120), .B1(n1281), .B2(n6689), .ZN(n6107) );
  OAI22_X2 U12885 ( .A1(n6688), .A2(n12120), .B1(n1187), .B2(n3689), .ZN(n6118) );
  INV_X4 U12886 ( .A(pipeline_csr_N674), .ZN(n12113) );
  OAI22_X2 U12887 ( .A1(n12255), .A2(n12118), .B1(n6821), .B2(n12113), .ZN(
        pipeline_csr_N1914) );
  OAI22_X2 U12888 ( .A1(n6703), .A2(n12120), .B1(n10544), .B2(n3683), .ZN(
        n6055) );
  INV_X4 U12889 ( .A(pipeline_csr_N770), .ZN(n12114) );
  OAI22_X2 U12890 ( .A1(n12615), .A2(n12118), .B1(n9403), .B2(n12114), .ZN(
        pipeline_csr_N2010) );
  INV_X4 U12891 ( .A(pipeline_csr_N706), .ZN(n12115) );
  OAI22_X2 U12892 ( .A1(n9469), .A2(n12118), .B1(n9404), .B2(n12115), .ZN(
        pipeline_csr_N1946) );
  NAND2_X2 U12893 ( .A1(pipeline_csr_N834), .A2(n12350), .ZN(n12116) );
  OAI221_X2 U12894 ( .B1(n12120), .B2(n6704), .C1(n1441), .C2(n12352), .A(
        n12116), .ZN(n5988) );
  INV_X4 U12895 ( .A(pipeline_csr_N738), .ZN(n12117) );
  OAI22_X2 U12896 ( .A1(n12612), .A2(n12118), .B1(n9406), .B2(n12117), .ZN(
        pipeline_csr_N1978) );
  NAND2_X2 U12897 ( .A1(pipeline_csr_N802), .A2(n12346), .ZN(n12119) );
  OAI221_X2 U12898 ( .B1(n12120), .B2(n12347), .C1(n10546), .C2(n12349), .A(
        n12119), .ZN(n6020) );
  OAI22_X2 U12899 ( .A1(n7208), .A2(n6691), .B1(n460), .B2(n9523), .ZN(n6360)
         );
  INV_X4 U12900 ( .A(n12182), .ZN(n12363) );
  MUX2_X2 U12901 ( .A(n12355), .B(n12357), .S(n6633), .Z(n12121) );
  NAND2_X2 U12902 ( .A1(n12121), .A2(n12783), .ZN(n12125) );
  NOR2_X2 U12903 ( .A1(n9513), .A2(n12122), .ZN(n12123) );
  OAI22_X2 U12904 ( .A1(n12128), .A2(n12791), .B1(n12794), .B2(n12127), .ZN(
        n12139) );
  NAND4_X2 U12905 ( .A1(n12132), .A2(n12131), .A3(n12130), .A4(n12129), .ZN(
        n12136) );
  AOI221_X2 U12906 ( .B1(n9510), .B2(n12136), .C1(n9511), .C2(n12135), .A(
        n12134), .ZN(n12137) );
  NOR2_X2 U12907 ( .A1(n12376), .A2(n12137), .ZN(n12138) );
  MUX2_X2 U12908 ( .A(n12139), .B(n12138), .S(n12800), .Z(n12140) );
  AOI221_X2 U12909 ( .B1(pipeline_alu_N62), .B2(n6813), .C1(pipeline_alu_N256), 
        .C2(n6812), .A(n12140), .ZN(n12141) );
  NAND2_X2 U12910 ( .A1(n12142), .A2(n12141), .ZN(dmem_haddr[3]) );
  MUX2_X2 U12911 ( .A(pipeline_alu_out_WB[3]), .B(dmem_haddr[3]), .S(n9523), 
        .Z(n5841) );
  OAI22_X2 U12912 ( .A1(n1907), .A2(n12806), .B1(n6923), .B2(n9515), .ZN(
        n12143) );
  AOI221_X2 U12913 ( .B1(pipeline_alu_out_WB[3]), .B2(n12809), .C1(n6670), 
        .C2(n12144), .A(n12143), .ZN(n12145) );
  INV_X4 U12914 ( .A(n12145), .ZN(n5809) );
  INV_X4 U12915 ( .A(pipeline_csr_N651), .ZN(n12146) );
  OAI22_X2 U12916 ( .A1(n12255), .A2(n12147), .B1(n6821), .B2(n12146), .ZN(
        pipeline_csr_N1891) );
  NAND3_X2 U12917 ( .A1(n6748), .A2(n13130), .A3(n7051), .ZN(n12621) );
  INV_X4 U12918 ( .A(n12150), .ZN(n12388) );
  NAND2_X2 U12919 ( .A1(pipeline_ctrl_prev_ex_code_WB[3]), .A2(n7215), .ZN(
        n12151) );
  OAI221_X2 U12920 ( .B1(n1482), .B2(n12620), .C1(n1907), .C2(n12621), .A(
        n12151), .ZN(n5972) );
  NAND2_X2 U12921 ( .A1(pipeline_csr_N304), .A2(n6750), .ZN(n12152) );
  OAI221_X2 U12922 ( .B1(n1486), .B2(n6687), .C1(n1907), .C2(n6705), .A(n12152), .ZN(n5872) );
  OAI22_X2 U12923 ( .A1(n1518), .A2(n6660), .B1(n1907), .B2(n9516), .ZN(n6210)
         );
  INV_X4 U12924 ( .A(n12622), .ZN(n1915) );
  INV_X4 U12925 ( .A(n12816), .ZN(n12153) );
  NAND2_X2 U12926 ( .A1(n12153), .A2(pipeline_csr_priv_stack_0), .ZN(n12154)
         );
  OAI221_X2 U12927 ( .B1(n12155), .B2(n12822), .C1(n1915), .C2(n12820), .A(
        n12154), .ZN(n6297) );
  INV_X4 U12928 ( .A(n12822), .ZN(n12157) );
  NOR2_X2 U12929 ( .A1(n12155), .A2(n12816), .ZN(n12156) );
  NOR2_X2 U12930 ( .A1(n12157), .A2(n12156), .ZN(n12158) );
  OAI221_X2 U12931 ( .B1(n1549), .B2(n12159), .C1(n1907), .C2(n12820), .A(
        n12158), .ZN(n5982) );
  OAI22_X2 U12932 ( .A1(n6701), .A2(n6691), .B1(n414), .B2(n9524), .ZN(n6337)
         );
  INV_X4 U12933 ( .A(n12160), .ZN(n12173) );
  NAND2_X2 U12934 ( .A1(n12161), .A2(n9511), .ZN(n12162) );
  NOR2_X2 U12935 ( .A1(n9513), .A2(n12166), .ZN(n12167) );
  OAI221_X2 U12936 ( .B1(n12169), .B2(n12168), .C1(n6601), .C2(n12167), .A(
        n12659), .ZN(n12170) );
  AOI221_X2 U12937 ( .B1(n12174), .B2(n12173), .C1(n12172), .C2(n12171), .A(
        n12170), .ZN(n12185) );
  MUX2_X2 U12938 ( .A(n12355), .B(n12357), .S(n6601), .Z(n12179) );
  NAND2_X2 U12939 ( .A1(n12179), .A2(n9512), .ZN(n12180) );
  OAI221_X2 U12940 ( .B1(n6746), .B2(n12639), .C1(n6811), .C2(n12182), .A(
        n12181), .ZN(n12183) );
  AOI221_X2 U12941 ( .B1(pipeline_alu_N86), .B2(n6813), .C1(pipeline_alu_N280), 
        .C2(n6812), .A(n12183), .ZN(n12184) );
  NAND2_X2 U12942 ( .A1(n12185), .A2(n12184), .ZN(dmem_haddr[27]) );
  MUX2_X2 U12943 ( .A(pipeline_alu_out_WB[27]), .B(dmem_haddr[27]), .S(n9524), 
        .Z(n5817) );
  OAI22_X2 U12944 ( .A1(n12805), .A2(n12186), .B1(n562), .B2(n9498), .ZN(
        n12187) );
  AOI221_X2 U12945 ( .B1(n12668), .B2(n12188), .C1(pipeline_alu_out_WB[27]), 
        .C2(n12809), .A(n12187), .ZN(n12189) );
  INV_X4 U12946 ( .A(n12189), .ZN(n5785) );
  NAND2_X2 U12947 ( .A1(pipeline_csr_N328), .A2(n6750), .ZN(n12190) );
  OAI221_X2 U12948 ( .B1(n12198), .B2(n6705), .C1(n1510), .C2(n6687), .A(
        n12190), .ZN(n5848) );
  OAI22_X2 U12949 ( .A1(n6659), .A2(n12198), .B1(n1282), .B2(n6689), .ZN(n6108) );
  OAI22_X2 U12950 ( .A1(n6688), .A2(n12198), .B1(n1188), .B2(n3689), .ZN(n6117) );
  INV_X4 U12951 ( .A(pipeline_csr_N675), .ZN(n12191) );
  OAI22_X2 U12952 ( .A1(n12255), .A2(n12196), .B1(n6821), .B2(n12191), .ZN(
        pipeline_csr_N1915) );
  OAI22_X2 U12953 ( .A1(n6703), .A2(n12198), .B1(n10468), .B2(n3683), .ZN(
        n6054) );
  INV_X4 U12954 ( .A(pipeline_csr_N771), .ZN(n12192) );
  OAI22_X2 U12955 ( .A1(n12615), .A2(n12196), .B1(n9403), .B2(n12192), .ZN(
        pipeline_csr_N2011) );
  INV_X4 U12956 ( .A(pipeline_csr_N707), .ZN(n12193) );
  OAI22_X2 U12957 ( .A1(n9469), .A2(n12196), .B1(n9404), .B2(n12193), .ZN(
        pipeline_csr_N1947) );
  NAND2_X2 U12958 ( .A1(pipeline_csr_N835), .A2(n12350), .ZN(n12194) );
  OAI221_X2 U12959 ( .B1(n12198), .B2(n6704), .C1(n1442), .C2(n12352), .A(
        n12194), .ZN(n5987) );
  INV_X4 U12960 ( .A(pipeline_csr_N739), .ZN(n12195) );
  OAI22_X2 U12961 ( .A1(n12612), .A2(n12196), .B1(n9406), .B2(n12195), .ZN(
        pipeline_csr_N1979) );
  NAND2_X2 U12962 ( .A1(pipeline_csr_N803), .A2(n12346), .ZN(n12197) );
  OAI221_X2 U12963 ( .B1(n12198), .B2(n12347), .C1(n10470), .C2(n12349), .A(
        n12197), .ZN(n6019) );
  OAI22_X2 U12964 ( .A1(n7209), .A2(n6691), .B1(n462), .B2(n9525), .ZN(n6361)
         );
  NAND2_X2 U12965 ( .A1(n9510), .A2(n12800), .ZN(n12577) );
  INV_X4 U12966 ( .A(n12577), .ZN(n12656) );
  NAND2_X2 U12967 ( .A1(n12656), .A2(n12199), .ZN(n12564) );
  INV_X4 U12968 ( .A(n12564), .ZN(n12643) );
  MUX2_X2 U12969 ( .A(n12355), .B(n12357), .S(n12200), .Z(n12201) );
  NAND2_X2 U12970 ( .A1(n12201), .A2(n12783), .ZN(n12207) );
  NAND2_X2 U12971 ( .A1(n9479), .A2(n12202), .ZN(n12203) );
  NAND2_X2 U12972 ( .A1(n12203), .A2(n12783), .ZN(n12204) );
  NAND2_X2 U12973 ( .A1(n12204), .A2(n6564), .ZN(n12205) );
  NAND2_X2 U12974 ( .A1(n12205), .A2(n12659), .ZN(n12206) );
  AOI221_X2 U12975 ( .B1(n12643), .B2(n12208), .C1(n12207), .C2(
        pipeline_alu_src_b[28]), .A(n12206), .ZN(n12231) );
  INV_X4 U12976 ( .A(n12209), .ZN(n12216) );
  INV_X4 U12977 ( .A(n12210), .ZN(n12215) );
  INV_X4 U12978 ( .A(n12211), .ZN(n12214) );
  INV_X4 U12979 ( .A(n12212), .ZN(n12213) );
  NOR4_X2 U12980 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12217) );
  NOR2_X2 U12981 ( .A1(n12217), .A2(n12577), .ZN(n12225) );
  INV_X4 U12982 ( .A(n12218), .ZN(n12223) );
  NAND2_X2 U12983 ( .A1(n9511), .A2(n12219), .ZN(n12220) );
  MUX2_X2 U12984 ( .A(n12223), .B(n12222), .S(n12800), .Z(n12224) );
  NOR2_X2 U12985 ( .A1(n12225), .A2(n12224), .ZN(n12228) );
  INV_X4 U12986 ( .A(n12226), .ZN(n12227) );
  OAI22_X2 U12987 ( .A1(n12228), .A2(n12590), .B1(n12227), .B2(n12639), .ZN(
        n12229) );
  AOI221_X2 U12988 ( .B1(pipeline_alu_N87), .B2(n6813), .C1(pipeline_alu_N281), 
        .C2(n6812), .A(n12229), .ZN(n12230) );
  NAND2_X2 U12989 ( .A1(n12231), .A2(n12230), .ZN(dmem_haddr[28]) );
  MUX2_X2 U12990 ( .A(pipeline_alu_out_WB[28]), .B(dmem_haddr[28]), .S(n9522), 
        .Z(n5816) );
  OAI22_X2 U12991 ( .A1(n12805), .A2(n12232), .B1(n563), .B2(n9498), .ZN(
        n12233) );
  AOI221_X2 U12992 ( .B1(n12668), .B2(n12234), .C1(pipeline_alu_out_WB[28]), 
        .C2(n12809), .A(n12233), .ZN(n12235) );
  INV_X4 U12993 ( .A(n12235), .ZN(n5784) );
  NAND2_X2 U12994 ( .A1(pipeline_csr_N329), .A2(n6750), .ZN(n12236) );
  OAI221_X2 U12995 ( .B1(n1511), .B2(n6687), .C1(n12242), .C2(n6705), .A(
        n12236), .ZN(n5847) );
  OAI22_X2 U12996 ( .A1(n6659), .A2(n12242), .B1(n1283), .B2(n6689), .ZN(n6109) );
  OAI22_X2 U12997 ( .A1(n6702), .A2(n12242), .B1(n10430), .B2(n9529), .ZN(
        n6148) );
  OAI22_X2 U12998 ( .A1(n6688), .A2(n12242), .B1(n1189), .B2(n3689), .ZN(n6116) );
  OAI22_X2 U12999 ( .A1(n6703), .A2(n12242), .B1(n1251), .B2(n3683), .ZN(n6053) );
  INV_X4 U13000 ( .A(pipeline_csr_N676), .ZN(n12237) );
  OAI22_X2 U13001 ( .A1(n12255), .A2(n12244), .B1(n6821), .B2(n12237), .ZN(
        pipeline_csr_N1916) );
  INV_X4 U13002 ( .A(pipeline_csr_N772), .ZN(n12238) );
  OAI22_X2 U13003 ( .A1(n12615), .A2(n12244), .B1(n9403), .B2(n12238), .ZN(
        pipeline_csr_N2012) );
  NAND2_X2 U13004 ( .A1(pipeline_csr_N836), .A2(n9476), .ZN(n12239) );
  OAI221_X2 U13005 ( .B1(n12242), .B2(n6704), .C1(n1443), .C2(n12352), .A(
        n12239), .ZN(n5986) );
  INV_X4 U13006 ( .A(pipeline_csr_N740), .ZN(n12240) );
  OAI22_X2 U13007 ( .A1(n12612), .A2(n12244), .B1(n9405), .B2(n12240), .ZN(
        pipeline_csr_N1980) );
  NAND2_X2 U13008 ( .A1(pipeline_csr_N804), .A2(n9472), .ZN(n12241) );
  OAI221_X2 U13009 ( .B1(n12242), .B2(n12347), .C1(n10433), .C2(n12349), .A(
        n12241), .ZN(n6018) );
  INV_X4 U13010 ( .A(pipeline_csr_N708), .ZN(n12243) );
  OAI22_X2 U13011 ( .A1(n9469), .A2(n12244), .B1(n12257), .B2(n12243), .ZN(
        pipeline_csr_N1948) );
  INV_X4 U13012 ( .A(pipeline_csr_N684), .ZN(n12245) );
  OAI22_X2 U13013 ( .A1(n9469), .A2(n12610), .B1(n9404), .B2(n12245), .ZN(
        pipeline_csr_N1924) );
  INV_X4 U13014 ( .A(pipeline_csr_N681), .ZN(n12246) );
  OAI22_X2 U13015 ( .A1(n9469), .A2(n12354), .B1(n12257), .B2(n12246), .ZN(
        pipeline_csr_N1921) );
  INV_X4 U13016 ( .A(pipeline_csr_N680), .ZN(n12247) );
  OAI22_X2 U13017 ( .A1(n12614), .A2(n9469), .B1(n12257), .B2(n12247), .ZN(
        pipeline_csr_N1920) );
  INV_X4 U13018 ( .A(pipeline_csr_N679), .ZN(n12248) );
  OAI22_X2 U13019 ( .A1(n6821), .A2(n12248), .B1(n12603), .B2(n12255), .ZN(
        pipeline_csr_N1919) );
  INV_X4 U13020 ( .A(pipeline_csr_N678), .ZN(n12249) );
  OAI22_X2 U13021 ( .A1(n6821), .A2(n12249), .B1(n12607), .B2(n12255), .ZN(
        pipeline_csr_N1918) );
  INV_X4 U13022 ( .A(pipeline_csr_N677), .ZN(n12250) );
  OAI22_X2 U13023 ( .A1(n12335), .A2(n12255), .B1(n6821), .B2(n12250), .ZN(
        pipeline_csr_N1917) );
  INV_X4 U13024 ( .A(pipeline_csr_N652), .ZN(n12251) );
  OAI22_X2 U13025 ( .A1(n12610), .A2(n12255), .B1(n6821), .B2(n12251), .ZN(
        pipeline_csr_N1892) );
  INV_X4 U13026 ( .A(pipeline_csr_N650), .ZN(n12252) );
  OAI22_X2 U13027 ( .A1(n12260), .A2(n12255), .B1(n6821), .B2(n12252), .ZN(
        pipeline_csr_N1890) );
  INV_X4 U13028 ( .A(pipeline_csr_N649), .ZN(n12253) );
  OAI22_X2 U13029 ( .A1(n12354), .A2(n12255), .B1(n6821), .B2(n12253), .ZN(
        pipeline_csr_N1889) );
  INV_X4 U13030 ( .A(pipeline_csr_N648), .ZN(n12254) );
  OAI22_X2 U13031 ( .A1(n12614), .A2(n12255), .B1(n6821), .B2(n12254), .ZN(
        pipeline_csr_N1888) );
  INV_X4 U13032 ( .A(pipeline_csr_N682), .ZN(n12256) );
  OAI22_X2 U13033 ( .A1(n9469), .A2(n12260), .B1(n9404), .B2(n12256), .ZN(
        pipeline_csr_N1922) );
  INV_X4 U13034 ( .A(pipeline_csr_N714), .ZN(n12259) );
  OAI22_X2 U13035 ( .A1(n12612), .A2(n12260), .B1(n9406), .B2(n12259), .ZN(
        pipeline_csr_N1954) );
  NAND2_X2 U13036 ( .A1(pipeline_csr_N778), .A2(n9472), .ZN(n12261) );
  OAI221_X2 U13037 ( .B1(n1909), .B2(n12347), .C1(n1385), .C2(n12349), .A(
        n12261), .ZN(n6044) );
  MUX2_X2 U13038 ( .A(n12355), .B(n12357), .S(n9399), .Z(n12262) );
  NAND2_X2 U13039 ( .A1(n12262), .A2(n12783), .ZN(n12267) );
  NOR2_X2 U13040 ( .A1(n9513), .A2(n12263), .ZN(n12264) );
  NOR2_X2 U13041 ( .A1(n9399), .A2(n12264), .ZN(n12266) );
  INV_X4 U13042 ( .A(n12269), .ZN(n12270) );
  OAI22_X2 U13043 ( .A1(n12271), .A2(n12791), .B1(n12794), .B2(n12270), .ZN(
        n12284) );
  INV_X4 U13044 ( .A(n12272), .ZN(n12280) );
  OAI22_X2 U13045 ( .A1(n12278), .A2(n12645), .B1(n12277), .B2(n9509), .ZN(
        n12279) );
  AOI221_X2 U13046 ( .B1(n12780), .B2(n12281), .C1(n9508), .C2(n12280), .A(
        n12279), .ZN(n12282) );
  NOR2_X2 U13047 ( .A1(n12376), .A2(n12282), .ZN(n12283) );
  MUX2_X2 U13048 ( .A(n12284), .B(n12283), .S(n12800), .Z(n12285) );
  AOI221_X2 U13049 ( .B1(pipeline_alu_N61), .B2(n6813), .C1(pipeline_alu_N255), 
        .C2(n6812), .A(n12285), .ZN(n12286) );
  NAND2_X2 U13050 ( .A1(n12287), .A2(n12286), .ZN(dmem_haddr[2]) );
  MUX2_X2 U13051 ( .A(pipeline_alu_out_WB[2]), .B(dmem_haddr[2]), .S(n9525), 
        .Z(n5842) );
  OAI22_X2 U13052 ( .A1(n1909), .A2(n12806), .B1(n9515), .B2(n12288), .ZN(
        n12289) );
  AOI221_X2 U13053 ( .B1(pipeline_alu_out_WB[2]), .B2(n12809), .C1(n6670), 
        .C2(n12290), .A(n12289), .ZN(n12291) );
  INV_X4 U13054 ( .A(n12291), .ZN(n5810) );
  NAND2_X2 U13055 ( .A1(n12388), .A2(n12292), .ZN(n12293) );
  OAI221_X2 U13056 ( .B1(n1481), .B2(n12620), .C1(n1909), .C2(n12621), .A(
        n12293), .ZN(n5973) );
  NAND2_X2 U13057 ( .A1(pipeline_csr_N303), .A2(n6750), .ZN(n12294) );
  OAI221_X2 U13058 ( .B1(n1485), .B2(n6687), .C1(n1909), .C2(n6705), .A(n12294), .ZN(n5873) );
  OAI22_X2 U13059 ( .A1(n1517), .A2(n6660), .B1(n1909), .B2(n9516), .ZN(n6209)
         );
  INV_X4 U13060 ( .A(n12295), .ZN(n12296) );
  OAI22_X2 U13061 ( .A1(n12296), .A2(n6691), .B1(n412), .B2(n9523), .ZN(n6336)
         );
  MUX2_X2 U13062 ( .A(n12355), .B(n12357), .S(n12297), .Z(n12298) );
  NAND2_X2 U13063 ( .A1(n12298), .A2(n12783), .ZN(n12304) );
  NAND2_X2 U13064 ( .A1(n9479), .A2(n12299), .ZN(n12300) );
  NAND2_X2 U13065 ( .A1(n12300), .A2(n12783), .ZN(n12301) );
  NAND2_X2 U13066 ( .A1(n12301), .A2(pipeline_alu_src_a[29]), .ZN(n12302) );
  NAND2_X2 U13067 ( .A1(n12302), .A2(n12659), .ZN(n12303) );
  AOI221_X2 U13068 ( .B1(n12305), .B2(n12643), .C1(n12304), .C2(n6556), .A(
        n12303), .ZN(n12327) );
  INV_X4 U13069 ( .A(n12306), .ZN(n12313) );
  INV_X4 U13070 ( .A(n12307), .ZN(n12312) );
  INV_X4 U13071 ( .A(n12308), .ZN(n12311) );
  INV_X4 U13072 ( .A(n12309), .ZN(n12310) );
  NOR4_X2 U13073 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12314) );
  NOR2_X2 U13074 ( .A1(n12314), .A2(n12577), .ZN(n12321) );
  NAND2_X2 U13075 ( .A1(n9511), .A2(n12315), .ZN(n12316) );
  MUX2_X2 U13076 ( .A(n12319), .B(n12318), .S(n12800), .Z(n12320) );
  NOR2_X2 U13077 ( .A1(n12321), .A2(n12320), .ZN(n12324) );
  INV_X4 U13078 ( .A(n12322), .ZN(n12323) );
  OAI22_X2 U13079 ( .A1(n12324), .A2(n12590), .B1(n12323), .B2(n12639), .ZN(
        n12325) );
  AOI221_X2 U13080 ( .B1(pipeline_alu_N88), .B2(n6813), .C1(pipeline_alu_N282), 
        .C2(n6812), .A(n12325), .ZN(n12326) );
  NAND2_X2 U13081 ( .A1(n12327), .A2(n12326), .ZN(dmem_haddr[29]) );
  MUX2_X2 U13082 ( .A(pipeline_alu_out_WB[29]), .B(dmem_haddr[29]), .S(n9522), 
        .Z(n5815) );
  OAI22_X2 U13083 ( .A1(n12805), .A2(n12328), .B1(n564), .B2(n9498), .ZN(
        n12329) );
  AOI221_X2 U13084 ( .B1(n12668), .B2(n12330), .C1(pipeline_alu_out_WB[29]), 
        .C2(n12809), .A(n12329), .ZN(n12331) );
  INV_X4 U13085 ( .A(n12331), .ZN(n5783) );
  NAND2_X2 U13086 ( .A1(pipeline_csr_N330), .A2(n6750), .ZN(n12332) );
  OAI221_X2 U13087 ( .B1(n12338), .B2(n6705), .C1(n1512), .C2(n6687), .A(
        n12332), .ZN(n5846) );
  OAI22_X2 U13088 ( .A1(n6659), .A2(n12338), .B1(n1284), .B2(n6689), .ZN(n6110) );
  OAI22_X2 U13089 ( .A1(n6702), .A2(n12338), .B1(n10362), .B2(n9529), .ZN(
        n6147) );
  OAI22_X2 U13090 ( .A1(n6688), .A2(n12338), .B1(n1190), .B2(n3689), .ZN(n6115) );
  OAI22_X2 U13091 ( .A1(n6703), .A2(n12338), .B1(n10365), .B2(n3683), .ZN(
        n6052) );
  INV_X4 U13092 ( .A(pipeline_csr_N773), .ZN(n12333) );
  OAI22_X2 U13093 ( .A1(n9492), .A2(n12335), .B1(n9403), .B2(n12333), .ZN(
        pipeline_csr_N2013) );
  NAND2_X2 U13094 ( .A1(pipeline_csr_N805), .A2(n9472), .ZN(n12334) );
  OAI221_X2 U13095 ( .B1(n12338), .B2(n12347), .C1(n10367), .C2(n12349), .A(
        n12334), .ZN(n6017) );
  INV_X4 U13096 ( .A(pipeline_csr_N741), .ZN(n12336) );
  OAI22_X2 U13097 ( .A1(n9406), .A2(n12336), .B1(n12612), .B2(n12335), .ZN(
        pipeline_csr_N1981) );
  NAND2_X2 U13098 ( .A1(pipeline_csr_N837), .A2(n9476), .ZN(n12337) );
  OAI221_X2 U13099 ( .B1(n12338), .B2(n6704), .C1(n1444), .C2(n12352), .A(
        n12337), .ZN(n6047) );
  INV_X4 U13100 ( .A(n12339), .ZN(n1905) );
  NAND2_X2 U13101 ( .A1(pipeline_csr_N812), .A2(n12350), .ZN(n12340) );
  OAI221_X2 U13102 ( .B1(n1905), .B2(n6704), .C1(n11231), .C2(n12352), .A(
        n12340), .ZN(n6010) );
  NAND2_X2 U13103 ( .A1(pipeline_csr_N808), .A2(n12350), .ZN(n12341) );
  OAI221_X2 U13104 ( .B1(n1915), .B2(n6704), .C1(n11259), .C2(n12352), .A(
        n12341), .ZN(n6014) );
  NAND2_X2 U13105 ( .A1(pipeline_csr_N807), .A2(n9472), .ZN(n12342) );
  OAI221_X2 U13106 ( .B1(n12601), .B2(n12347), .C1(n10293), .C2(n12349), .A(
        n12342), .ZN(n6015) );
  NAND2_X2 U13107 ( .A1(pipeline_csr_N806), .A2(n9472), .ZN(n12343) );
  OAI221_X2 U13108 ( .B1(n12670), .B2(n12347), .C1(n10252), .C2(n12349), .A(
        n12343), .ZN(n6016) );
  NAND2_X2 U13109 ( .A1(pipeline_csr_N780), .A2(n9472), .ZN(n12344) );
  OAI221_X2 U13110 ( .B1(n1905), .B2(n12347), .C1(n1387), .C2(n12349), .A(
        n12344), .ZN(n6042) );
  NAND2_X2 U13111 ( .A1(pipeline_csr_N777), .A2(n9472), .ZN(n12345) );
  OAI221_X2 U13112 ( .B1(n1911), .B2(n12347), .C1(n1384), .C2(n12349), .A(
        n12345), .ZN(n6045) );
  NAND2_X2 U13113 ( .A1(n9474), .A2(n12622), .ZN(n12348) );
  OAI221_X2 U13114 ( .B1(pipeline_csr_instret_full[0]), .B2(n9473), .C1(n1319), 
        .C2(n12349), .A(n12348), .ZN(n6046) );
  NAND2_X2 U13115 ( .A1(pipeline_csr_N809), .A2(n12350), .ZN(n12351) );
  OAI221_X2 U13116 ( .B1(n1911), .B2(n6704), .C1(n10317), .C2(n12352), .A(
        n12351), .ZN(n6013) );
  INV_X4 U13117 ( .A(pipeline_csr_N713), .ZN(n12353) );
  OAI22_X2 U13118 ( .A1(n12612), .A2(n12354), .B1(n9405), .B2(n12353), .ZN(
        pipeline_csr_N1953) );
  MUX2_X2 U13119 ( .A(n12355), .B(n12357), .S(n6631), .Z(n12356) );
  NAND2_X2 U13120 ( .A1(n12356), .A2(n12783), .ZN(n12361) );
  NOR2_X2 U13121 ( .A1(n9513), .A2(n12358), .ZN(n12359) );
  INV_X4 U13122 ( .A(n12364), .ZN(n12365) );
  OAI22_X2 U13123 ( .A1(n12366), .A2(n12791), .B1(n12794), .B2(n12365), .ZN(
        n12378) );
  NAND2_X2 U13124 ( .A1(n9489), .A2(n6632), .ZN(n12368) );
  NAND4_X2 U13125 ( .A1(n12370), .A2(n12369), .A3(n12368), .A4(n12367), .ZN(
        n12374) );
  OAI22_X2 U13126 ( .A1(n6801), .A2(n9507), .B1(n12371), .B2(n12582), .ZN(
        n12372) );
  AOI221_X2 U13127 ( .B1(n9510), .B2(n12374), .C1(n9511), .C2(n12373), .A(
        n12372), .ZN(n12375) );
  NOR2_X2 U13128 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  MUX2_X2 U13129 ( .A(n12378), .B(n12377), .S(n12800), .Z(n12379) );
  AOI221_X2 U13130 ( .B1(pipeline_alu_N60), .B2(n6813), .C1(pipeline_alu_N254), 
        .C2(n6812), .A(n12379), .ZN(n12380) );
  NAND2_X2 U13131 ( .A1(n12381), .A2(n12380), .ZN(dmem_haddr[1]) );
  MUX2_X2 U13132 ( .A(pipeline_alu_out_WB[1]), .B(dmem_haddr[1]), .S(n9524), 
        .Z(n5843) );
  INV_X4 U13133 ( .A(imem_haddr[1]), .ZN(n12382) );
  OAI22_X2 U13134 ( .A1(n12535), .A2(n9494), .B1(n9493), .B2(n12382), .ZN(
        n5970) );
  OAI22_X2 U13135 ( .A1(n12535), .A2(n9496), .B1(n716), .B2(n6662), .ZN(n5937)
         );
  MUX2_X2 U13136 ( .A(n12383), .B(pipeline_PC_DX[1]), .S(n9523), .Z(n5936) );
  OAI22_X2 U13137 ( .A1(n536), .A2(n9498), .B1(n12936), .B2(n12617), .ZN(
        n12384) );
  AOI221_X2 U13138 ( .B1(pipeline_csr_mbadaddr[1]), .B2(n9514), .C1(n12668), 
        .C2(n12385), .A(n12384), .ZN(n12386) );
  INV_X4 U13139 ( .A(n12386), .ZN(n5811) );
  NOR2_X2 U13140 ( .A1(pipeline_ctrl_wr_reg_unkilled_WB), .A2(
        pipeline_ctrl_had_ex_WB), .ZN(n12389) );
  OAI22_X2 U13141 ( .A1(n1911), .A2(n12621), .B1(n1480), .B2(n12620), .ZN(
        n12387) );
  AOI221_X2 U13142 ( .B1(n12389), .B2(n12388), .C1(n7215), .C2(
        pipeline_ctrl_prev_ex_code_WB[1]), .A(n12387), .ZN(n12390) );
  INV_X4 U13143 ( .A(n12390), .ZN(n5974) );
  NOR2_X2 U13144 ( .A1(n1484), .A2(n6687), .ZN(n5874) );
  OAI22_X2 U13145 ( .A1(n1516), .A2(n6660), .B1(n1911), .B2(n9516), .ZN(n6208)
         );
  INV_X4 U13146 ( .A(n12391), .ZN(n12392) );
  OAI22_X2 U13147 ( .A1(n12392), .A2(n6691), .B1(n410), .B2(n9525), .ZN(n6335)
         );
  OAI22_X2 U13148 ( .A1(n1905), .A2(n6690), .B1(n1195), .B2(n6708), .ZN(n6204)
         );
  NAND2_X2 U13149 ( .A1(pipeline_csr_N332), .A2(n6750), .ZN(n12393) );
  OAI221_X2 U13150 ( .B1(n1514), .B2(n6687), .C1(n12601), .C2(n6705), .A(
        n12393), .ZN(n5844) );
  NAND3_X2 U13151 ( .A1(n12406), .A2(n6799), .A3(n12396), .ZN(n12560) );
  INV_X4 U13152 ( .A(n12560), .ZN(n12409) );
  NAND3_X2 U13153 ( .A1(n13097), .A2(n12397), .A3(n12409), .ZN(n12404) );
  INV_X4 U13154 ( .A(n12398), .ZN(n12400) );
  NAND2_X2 U13155 ( .A1(n12400), .A2(n12399), .ZN(n12401) );
  NAND4_X2 U13156 ( .A1(n12406), .A2(n12402), .A3(n13097), .A4(n12401), .ZN(
        n12403) );
  NAND2_X2 U13157 ( .A1(n12406), .A2(n12405), .ZN(n12407) );
  INV_X4 U13158 ( .A(n12407), .ZN(n12412) );
  AOI221_X2 U13159 ( .B1(pipeline_PC_DX[31]), .B2(n9337), .C1(
        pipeline_handler_PC[31]), .C2(n6630), .A(n12414), .ZN(n12415) );
  OAI221_X2 U13160 ( .B1(n9487), .B2(n12416), .C1(n1514), .C2(n6661), .A(
        n12415), .ZN(pipeline_PCmux_base[31]) );
  NAND2_X2 U13161 ( .A1(pipeline_csr_N331), .A2(n6750), .ZN(n12417) );
  OAI221_X2 U13162 ( .B1(n12670), .B2(n6705), .C1(n1513), .C2(n6687), .A(
        n12417), .ZN(n5845) );
  NOR2_X2 U13163 ( .A1(n12418), .A2(n9484), .ZN(n12419) );
  AOI221_X2 U13164 ( .B1(pipeline_PC_DX[30]), .B2(n9480), .C1(
        pipeline_handler_PC[30]), .C2(n6630), .A(n12419), .ZN(n12420) );
  OAI221_X2 U13165 ( .B1(n9488), .B2(n12421), .C1(n1513), .C2(n6661), .A(
        n12420), .ZN(pipeline_PCmux_base[30]) );
  AOI221_X2 U13166 ( .B1(pipeline_PC_DX[29]), .B2(n9480), .C1(
        pipeline_handler_PC[29]), .C2(n6630), .A(n12423), .ZN(n12424) );
  OAI221_X2 U13167 ( .B1(n9488), .B2(n12425), .C1(n1512), .C2(n6661), .A(
        n12424), .ZN(pipeline_PCmux_base[29]) );
  AOI221_X2 U13168 ( .B1(pipeline_PC_DX[27]), .B2(n9482), .C1(
        pipeline_handler_PC[27]), .C2(n6630), .A(n12431), .ZN(n12432) );
  OAI221_X2 U13169 ( .B1(n9488), .B2(n12433), .C1(n1510), .C2(n6661), .A(
        n12432), .ZN(pipeline_PCmux_base[27]) );
  NOR2_X2 U13170 ( .A1(n12434), .A2(n9484), .ZN(n12435) );
  AOI221_X2 U13171 ( .B1(pipeline_PC_DX[26]), .B2(n6969), .C1(
        pipeline_handler_PC[26]), .C2(n6630), .A(n12435), .ZN(n12436) );
  OAI221_X2 U13172 ( .B1(n9488), .B2(n12437), .C1(n1509), .C2(n6661), .A(
        n12436), .ZN(pipeline_PCmux_base[26]) );
  NOR2_X2 U13173 ( .A1(n12438), .A2(n9484), .ZN(n12439) );
  AOI221_X2 U13174 ( .B1(pipeline_PC_DX[25]), .B2(n6969), .C1(
        pipeline_handler_PC[25]), .C2(n6630), .A(n12439), .ZN(n12440) );
  OAI221_X2 U13175 ( .B1(n9488), .B2(n12441), .C1(n1508), .C2(n6661), .A(
        n12440), .ZN(pipeline_PCmux_base[25]) );
  NOR2_X2 U13176 ( .A1(n12446), .A2(n9484), .ZN(n12447) );
  AOI221_X2 U13177 ( .B1(pipeline_PC_DX[23]), .B2(n6969), .C1(
        pipeline_handler_PC[23]), .C2(n6630), .A(n12447), .ZN(n12448) );
  OAI221_X2 U13178 ( .B1(n9488), .B2(n12449), .C1(n1506), .C2(n6661), .A(
        n12448), .ZN(pipeline_PCmux_base[23]) );
  NOR2_X2 U13179 ( .A1(n12450), .A2(n9484), .ZN(n12451) );
  AOI221_X2 U13180 ( .B1(pipeline_PC_DX[22]), .B2(n9480), .C1(
        pipeline_handler_PC[22]), .C2(n6630), .A(n12451), .ZN(n12452) );
  NOR2_X2 U13181 ( .A1(n12454), .A2(n9484), .ZN(n12455) );
  OAI221_X2 U13182 ( .B1(n9488), .B2(n12461), .C1(n1503), .C2(n6661), .A(
        n12460), .ZN(pipeline_PCmux_base[20]) );
  AOI221_X2 U13183 ( .B1(pipeline_PC_DX[19]), .B2(n6958), .C1(
        pipeline_handler_PC[19]), .C2(n6630), .A(n12463), .ZN(n12464) );
  NOR2_X2 U13184 ( .A1(n12466), .A2(n9485), .ZN(n12467) );
  AOI221_X2 U13185 ( .B1(pipeline_PC_DX[18]), .B2(n9480), .C1(
        pipeline_handler_PC[18]), .C2(n6630), .A(n12467), .ZN(n12468) );
  NOR2_X2 U13186 ( .A1(n12470), .A2(n9485), .ZN(n12471) );
  AOI221_X2 U13187 ( .B1(pipeline_PC_DX[17]), .B2(n6969), .C1(
        pipeline_handler_PC[17]), .C2(n6630), .A(n12471), .ZN(n12472) );
  OAI221_X2 U13188 ( .B1(n9488), .B2(n12480), .C1(n1498), .C2(n6661), .A(
        n12479), .ZN(pipeline_PCmux_base[15]) );
  AOI221_X2 U13189 ( .B1(pipeline_PC_DX[13]), .B2(n6958), .C1(
        pipeline_handler_PC[13]), .C2(n6630), .A(n12486), .ZN(n12487) );
  OAI221_X2 U13190 ( .B1(n9487), .B2(n12496), .C1(n1494), .C2(n6661), .A(
        n12495), .ZN(pipeline_PCmux_base[11]) );
  NOR2_X2 U13191 ( .A1(n12497), .A2(n9485), .ZN(n12498) );
  AOI221_X2 U13192 ( .B1(pipeline_PC_DX[10]), .B2(n9336), .C1(
        pipeline_handler_PC[10]), .C2(n6630), .A(n12498), .ZN(n12499) );
  OAI221_X2 U13193 ( .B1(n9487), .B2(n12500), .C1(n1493), .C2(n6661), .A(
        n12499), .ZN(pipeline_PCmux_base[10]) );
  AOI221_X2 U13194 ( .B1(n9337), .B2(pipeline_PC_DX[9]), .C1(
        pipeline_handler_PC[9]), .C2(n6630), .A(n12502), .ZN(n12503) );
  OAI221_X2 U13195 ( .B1(n9487), .B2(n12504), .C1(n1492), .C2(n6661), .A(
        n12503), .ZN(pipeline_PCmux_base[9]) );
  AOI221_X2 U13196 ( .B1(pipeline_PC_DX[8]), .B2(n6958), .C1(
        pipeline_handler_PC[8]), .C2(n6630), .A(n12506), .ZN(n12507) );
  OAI221_X2 U13197 ( .B1(n9487), .B2(n12508), .C1(n1491), .C2(n6661), .A(
        n12507), .ZN(pipeline_PCmux_base[8]) );
  AOI221_X2 U13198 ( .B1(pipeline_PC_DX[7]), .B2(n6958), .C1(
        pipeline_handler_PC[7]), .C2(n6630), .A(n12510), .ZN(n12511) );
  OAI221_X2 U13199 ( .B1(n9488), .B2(n12512), .C1(n1490), .C2(n6661), .A(
        n12511), .ZN(pipeline_PCmux_base[7]) );
  NOR2_X2 U13200 ( .A1(n12517), .A2(n9486), .ZN(n12518) );
  AOI221_X2 U13201 ( .B1(pipeline_PC_DX[5]), .B2(n9337), .C1(
        pipeline_handler_PC[5]), .C2(n6630), .A(n12518), .ZN(n12519) );
  OAI221_X2 U13202 ( .B1(n9487), .B2(n12520), .C1(n1488), .C2(n6661), .A(
        n12519), .ZN(pipeline_PCmux_base[5]) );
  NAND2_X2 U13203 ( .A1(pipeline_csr_N305), .A2(n6750), .ZN(n12521) );
  OAI221_X2 U13204 ( .B1(n1487), .B2(n6687), .C1(n1905), .C2(n6705), .A(n12521), .ZN(n5871) );
  OAI221_X2 U13205 ( .B1(n9487), .B2(n12525), .C1(n1487), .C2(n6661), .A(
        n12524), .ZN(pipeline_PCmux_base[4]) );
  AOI221_X2 U13206 ( .B1(pipeline_PC_DX[3]), .B2(n9336), .C1(
        pipeline_handler_PC[3]), .C2(n6630), .A(n12527), .ZN(n12528) );
  OAI221_X2 U13207 ( .B1(n9487), .B2(n12529), .C1(n1486), .C2(n6661), .A(
        n12528), .ZN(pipeline_PCmux_base[3]) );
  OAI22_X2 U13208 ( .A1(n1484), .A2(n6661), .B1(n9488), .B2(n12535), .ZN(
        n12536) );
  INV_X4 U13209 ( .A(n12537), .ZN(pipeline_PCmux_base[1]) );
  INV_X4 U13210 ( .A(imem_haddr[0]), .ZN(n12538) );
  OAI22_X2 U13211 ( .A1(n12539), .A2(n9494), .B1(n9493), .B2(n12538), .ZN(
        n5971) );
  OAI22_X2 U13212 ( .A1(n12539), .A2(n9496), .B1(n715), .B2(n6662), .ZN(n5939)
         );
  NOR2_X2 U13213 ( .A1(n1483), .A2(n6687), .ZN(n5875) );
  INV_X4 U13214 ( .A(n12541), .ZN(pipeline_PCmux_base[0]) );
  NAND2_X2 U13215 ( .A1(n12561), .A2(n9486), .ZN(n12543) );
  NAND2_X2 U13216 ( .A1(pipeline_imm_31_), .A2(n12543), .ZN(n12552) );
  INV_X4 U13217 ( .A(n12557), .ZN(n12550) );
  NAND2_X2 U13218 ( .A1(n12550), .A2(pipeline_regfile_N16), .ZN(n12544) );
  NAND2_X2 U13219 ( .A1(n12552), .A2(n12544), .ZN(pipeline_PCmux_offset[19])
         );
  NAND2_X2 U13220 ( .A1(n12550), .A2(pipeline_regfile_N15), .ZN(n12545) );
  NAND2_X2 U13221 ( .A1(n12552), .A2(n12545), .ZN(pipeline_PCmux_offset[18])
         );
  NAND2_X2 U13222 ( .A1(n12550), .A2(n12546), .ZN(n12547) );
  NAND2_X2 U13223 ( .A1(n12550), .A2(pipeline_dmem_type_2_), .ZN(n12548) );
  NAND2_X2 U13224 ( .A1(n12550), .A2(dmem_hsize[1]), .ZN(n12549) );
  NAND2_X2 U13225 ( .A1(n12550), .A2(dmem_hsize[0]), .ZN(n12551) );
  NOR2_X2 U13226 ( .A1(n713), .A2(n12555), .ZN(pipeline_PCmux_offset[10]) );
  NOR2_X2 U13227 ( .A1(n9632), .A2(n12555), .ZN(pipeline_PCmux_offset[9]) );
  NOR2_X2 U13228 ( .A1(n9634), .A2(n12555), .ZN(pipeline_PCmux_offset[8]) );
  NOR2_X2 U13229 ( .A1(n10236), .A2(n12555), .ZN(pipeline_PCmux_offset[7]) );
  NOR2_X2 U13230 ( .A1(n10338), .A2(n12555), .ZN(pipeline_PCmux_offset[6]) );
  NOR2_X2 U13231 ( .A1(n10336), .A2(n12555), .ZN(pipeline_PCmux_offset[5]) );
  NAND2_X2 U13232 ( .A1(n12557), .A2(n9486), .ZN(n12558) );
  INV_X4 U13233 ( .A(n12558), .ZN(n12562) );
  OAI22_X2 U13234 ( .A1(n8223), .A2(n12562), .B1(n597), .B2(n12561), .ZN(
        pipeline_PCmux_offset[3]) );
  NAND2_X2 U13235 ( .A1(n12558), .A2(pipeline_regfile_N19), .ZN(n12559) );
  OAI221_X2 U13236 ( .B1(n596), .B2(n12561), .C1(n12560), .C2(n9487), .A(
        n12559), .ZN(pipeline_PCmux_offset[2]) );
  OAI22_X2 U13237 ( .A1(n12416), .A2(n9494), .B1(n9493), .B2(n12563), .ZN(
        n5940) );
  OAI22_X2 U13238 ( .A1(n12416), .A2(n9497), .B1(n746), .B2(n6662), .ZN(n5877)
         );
  NOR2_X2 U13239 ( .A1(n12565), .A2(n12564), .ZN(n12569) );
  MUX2_X2 U13240 ( .A(n12793), .B(n9479), .S(n12566), .Z(n12568) );
  NOR4_X2 U13241 ( .A1(n12569), .A2(n12568), .A3(n9513), .A4(n12567), .ZN(
        n12592) );
  INV_X4 U13242 ( .A(n12570), .ZN(n12575) );
  INV_X4 U13243 ( .A(n12571), .ZN(n12574) );
  INV_X4 U13244 ( .A(n12572), .ZN(n12573) );
  NOR4_X2 U13245 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12578) );
  NOR2_X2 U13246 ( .A1(n12578), .A2(n12577), .ZN(n12586) );
  NAND2_X2 U13247 ( .A1(n9511), .A2(n12579), .ZN(n12580) );
  MUX2_X2 U13248 ( .A(n12584), .B(n12583), .S(n12800), .Z(n12585) );
  NOR2_X2 U13249 ( .A1(n12586), .A2(n12585), .ZN(n12591) );
  NAND2_X2 U13250 ( .A1(n9479), .A2(n12593), .ZN(n12587) );
  NAND2_X2 U13251 ( .A1(n12587), .A2(n12783), .ZN(n12588) );
  OAI221_X2 U13252 ( .B1(n12593), .B2(n12592), .C1(n12591), .C2(n12590), .A(
        n12589), .ZN(n12594) );
  MUX2_X2 U13253 ( .A(pipeline_alu_out_WB[31]), .B(dmem_haddr[31]), .S(n9524), 
        .Z(n5813) );
  OAI22_X2 U13254 ( .A1(n12601), .A2(n12806), .B1(n9515), .B2(n12595), .ZN(
        n12596) );
  AOI221_X2 U13255 ( .B1(pipeline_alu_out_WB[31]), .B2(n12809), .C1(n6670), 
        .C2(n12597), .A(n12596), .ZN(n12598) );
  INV_X4 U13256 ( .A(n12598), .ZN(n5781) );
  OAI221_X2 U13257 ( .B1(n1478), .B2(n12620), .C1(n12601), .C2(n12621), .A(
        n12624), .ZN(n5983) );
  OAI22_X2 U13258 ( .A1(n6659), .A2(n12601), .B1(n1286), .B2(n6689), .ZN(n6367) );
  OAI22_X2 U13259 ( .A1(n6702), .A2(n12601), .B1(n10287), .B2(n9529), .ZN(
        n6145) );
  OAI22_X2 U13260 ( .A1(n6688), .A2(n12601), .B1(n1192), .B2(n3689), .ZN(n6113) );
  OAI22_X2 U13261 ( .A1(n6703), .A2(n12601), .B1(n1254), .B2(n3683), .ZN(n6050) );
  INV_X4 U13262 ( .A(pipeline_csr_N743), .ZN(n12602) );
  OAI22_X2 U13263 ( .A1(n9405), .A2(n12602), .B1(n12612), .B2(n12603), .ZN(
        pipeline_csr_N1983) );
  INV_X4 U13264 ( .A(pipeline_csr_N775), .ZN(n12604) );
  OAI22_X2 U13265 ( .A1(n9403), .A2(n12604), .B1(n9492), .B2(n12603), .ZN(
        pipeline_csr_N2015) );
  INV_X4 U13266 ( .A(pipeline_csr_N774), .ZN(n12605) );
  OAI22_X2 U13267 ( .A1(n9403), .A2(n12605), .B1(n9492), .B2(n12607), .ZN(
        pipeline_csr_N2014) );
  INV_X4 U13268 ( .A(pipeline_csr_N748), .ZN(n12606) );
  OAI22_X2 U13269 ( .A1(n9492), .A2(n12610), .B1(n9403), .B2(n12606), .ZN(
        pipeline_csr_N1988) );
  INV_X4 U13270 ( .A(pipeline_csr_N742), .ZN(n12608) );
  OAI22_X2 U13271 ( .A1(n9406), .A2(n12608), .B1(n12612), .B2(n12607), .ZN(
        pipeline_csr_N1982) );
  INV_X4 U13272 ( .A(pipeline_csr_N716), .ZN(n12609) );
  OAI22_X2 U13273 ( .A1(n12612), .A2(n12610), .B1(n9405), .B2(n12609), .ZN(
        pipeline_csr_N1956) );
  INV_X4 U13274 ( .A(pipeline_csr_N712), .ZN(n12611) );
  OAI22_X2 U13275 ( .A1(n12614), .A2(n12612), .B1(n9406), .B2(n12611), .ZN(
        pipeline_csr_N1952) );
  INV_X4 U13276 ( .A(pipeline_csr_N744), .ZN(n12613) );
  OAI22_X2 U13277 ( .A1(n9492), .A2(n12614), .B1(n9403), .B2(n12613), .ZN(
        pipeline_csr_N1984) );
  MUX2_X2 U13278 ( .A(pipeline_alu_out_WB[0]), .B(dmem_haddr[0]), .S(n9525), 
        .Z(n6301) );
  MUX2_X2 U13279 ( .A(n12616), .B(pipeline_PC_DX[0]), .S(n9524), .Z(n5938) );
  OAI22_X2 U13280 ( .A1(n535), .A2(n9498), .B1(n12937), .B2(n12617), .ZN(
        n12618) );
  AOI221_X2 U13281 ( .B1(pipeline_csr_mbadaddr[0]), .B2(n9514), .C1(n12668), 
        .C2(n12622), .A(n12618), .ZN(n12619) );
  INV_X4 U13282 ( .A(n12619), .ZN(n5812) );
  INV_X4 U13283 ( .A(n12620), .ZN(n12628) );
  INV_X4 U13284 ( .A(n12621), .ZN(n12623) );
  NAND2_X2 U13285 ( .A1(n12623), .A2(n12622), .ZN(n12625) );
  NAND2_X2 U13286 ( .A1(n12625), .A2(n12624), .ZN(n12626) );
  AOI221_X2 U13287 ( .B1(pipeline_ctrl_prev_ex_code_WB[0]), .B2(n7215), .C1(
        n12628), .C2(n12627), .A(n12626), .ZN(n12629) );
  INV_X4 U13288 ( .A(n12629), .ZN(n5975) );
  OAI22_X2 U13289 ( .A1(n1515), .A2(n6660), .B1(n1915), .B2(n9516), .ZN(n6239)
         );
  INV_X4 U13290 ( .A(n12630), .ZN(n12631) );
  OAI22_X2 U13291 ( .A1(n12631), .A2(n6691), .B1(n408), .B2(n9524), .ZN(n6334)
         );
  OAI22_X2 U13292 ( .A1(n12421), .A2(n12632), .B1(n9493), .B2(n6953), .ZN(
        n5941) );
  OAI22_X2 U13293 ( .A1(n12421), .A2(n9497), .B1(n745), .B2(n6662), .ZN(n5879)
         );
  NAND2_X2 U13294 ( .A1(n9479), .A2(n12638), .ZN(n12633) );
  NAND2_X2 U13295 ( .A1(n12633), .A2(n12783), .ZN(n12644) );
  INV_X4 U13296 ( .A(n12634), .ZN(n12640) );
  MUX2_X2 U13297 ( .A(n12793), .B(n9479), .S(n12635), .Z(n12636) );
  NOR2_X2 U13298 ( .A1(n9513), .A2(n12636), .ZN(n12637) );
  OAI22_X2 U13299 ( .A1(n12640), .A2(n12639), .B1(n12638), .B2(n12637), .ZN(
        n12641) );
  AOI221_X2 U13300 ( .B1(n12644), .B2(n6997), .C1(n12643), .C2(n12642), .A(
        n12641), .ZN(n12664) );
  NOR2_X2 U13301 ( .A1(n6800), .A2(n12645), .ZN(n12646) );
  AOI221_X2 U13302 ( .B1(n9508), .B2(n12648), .C1(n12647), .C2(n12780), .A(
        n12646), .ZN(n12649) );
  MUX2_X2 U13303 ( .A(n12650), .B(n12649), .S(n12800), .Z(n12658) );
  NAND2_X2 U13304 ( .A1(n9489), .A2(n6997), .ZN(n12652) );
  NAND4_X2 U13305 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        n12655) );
  NAND2_X2 U13306 ( .A1(n12656), .A2(n12655), .ZN(n12657) );
  NAND2_X2 U13307 ( .A1(n12658), .A2(n12657), .ZN(n12661) );
  NAND2_X2 U13308 ( .A1(pipeline_alu_N283), .A2(n6812), .ZN(n12660) );
  MUX2_X2 U13309 ( .A(pipeline_alu_out_WB[30]), .B(dmem_haddr[30]), .S(n9525), 
        .Z(n5814) );
  OAI22_X2 U13310 ( .A1(n12805), .A2(n12665), .B1(n565), .B2(n9498), .ZN(
        n12666) );
  AOI221_X2 U13311 ( .B1(n12668), .B2(n12667), .C1(pipeline_alu_out_WB[30]), 
        .C2(n12809), .A(n12666), .ZN(n12669) );
  INV_X4 U13312 ( .A(n12669), .ZN(n5782) );
  OAI22_X2 U13313 ( .A1(n6659), .A2(n12670), .B1(n1285), .B2(n6689), .ZN(n6111) );
  OAI22_X2 U13314 ( .A1(n6702), .A2(n12670), .B1(n10243), .B2(n9529), .ZN(
        n6146) );
  OAI22_X2 U13315 ( .A1(n6688), .A2(n12670), .B1(n1191), .B2(n3689), .ZN(n6114) );
  OAI22_X2 U13316 ( .A1(n6703), .A2(n12670), .B1(n10249), .B2(n3683), .ZN(
        n6051) );
  OAI22_X2 U13317 ( .A1(n7211), .A2(n6691), .B1(n468), .B2(n9523), .ZN(n6364)
         );
  INV_X4 U13318 ( .A(pipeline_md_N281), .ZN(n12671) );
  OAI22_X2 U13319 ( .A1(n13058), .A2(n9504), .B1(n9505), .B2(n12671), .ZN(
        n12672) );
  AOI221_X2 U13320 ( .B1(pipeline_md_N59), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[30]), .A(n12672), .ZN(n12673) );
  INV_X4 U13321 ( .A(n12673), .ZN(n5683) );
  MUX2_X2 U13322 ( .A(pipeline_md_resp_result[30]), .B(pipeline_md_a[30]), .S(
        n9499), .Z(pipeline_md_result_muxed[30]) );
  MUX2_X2 U13323 ( .A(pipeline_md_resp_result[29]), .B(pipeline_md_a[29]), .S(
        n9499), .Z(pipeline_md_result_muxed[29]) );
  MUX2_X2 U13324 ( .A(pipeline_md_resp_result[28]), .B(pipeline_md_a[28]), .S(
        n9499), .Z(pipeline_md_result_muxed[28]) );
  MUX2_X2 U13325 ( .A(pipeline_md_resp_result[27]), .B(pipeline_md_a[27]), .S(
        n9499), .Z(pipeline_md_result_muxed[27]) );
  MUX2_X2 U13326 ( .A(pipeline_md_resp_result[26]), .B(pipeline_md_a[26]), .S(
        n9500), .Z(pipeline_md_result_muxed[26]) );
  MUX2_X2 U13327 ( .A(pipeline_md_resp_result[25]), .B(pipeline_md_a[25]), .S(
        n9499), .Z(pipeline_md_result_muxed[25]) );
  MUX2_X2 U13328 ( .A(pipeline_md_resp_result[24]), .B(pipeline_md_a[24]), .S(
        n9500), .Z(pipeline_md_result_muxed[24]) );
  MUX2_X2 U13329 ( .A(pipeline_md_resp_result[23]), .B(pipeline_md_a[23]), .S(
        n9500), .Z(pipeline_md_result_muxed[23]) );
  MUX2_X2 U13330 ( .A(pipeline_md_resp_result[22]), .B(pipeline_md_a[22]), .S(
        n9499), .Z(pipeline_md_result_muxed[22]) );
  MUX2_X2 U13331 ( .A(pipeline_md_resp_result[21]), .B(pipeline_md_a[21]), .S(
        n9500), .Z(pipeline_md_result_muxed[21]) );
  MUX2_X2 U13332 ( .A(pipeline_md_resp_result[20]), .B(pipeline_md_a[20]), .S(
        n9499), .Z(pipeline_md_result_muxed[20]) );
  MUX2_X2 U13333 ( .A(pipeline_md_resp_result[19]), .B(pipeline_md_a[19]), .S(
        n9500), .Z(pipeline_md_result_muxed[19]) );
  MUX2_X2 U13334 ( .A(pipeline_md_resp_result[18]), .B(pipeline_md_a[18]), .S(
        n9499), .Z(pipeline_md_result_muxed[18]) );
  MUX2_X2 U13335 ( .A(pipeline_md_resp_result[17]), .B(pipeline_md_a[17]), .S(
        n9500), .Z(pipeline_md_result_muxed[17]) );
  MUX2_X2 U13336 ( .A(pipeline_md_resp_result[16]), .B(pipeline_md_a[16]), .S(
        n9500), .Z(pipeline_md_result_muxed[16]) );
  MUX2_X2 U13337 ( .A(pipeline_md_resp_result[15]), .B(pipeline_md_a[15]), .S(
        n9499), .Z(pipeline_md_result_muxed[15]) );
  MUX2_X2 U13338 ( .A(pipeline_md_resp_result[14]), .B(pipeline_md_a[14]), .S(
        n9500), .Z(pipeline_md_result_muxed[14]) );
  MUX2_X2 U13339 ( .A(pipeline_md_resp_result[13]), .B(pipeline_md_a[13]), .S(
        n9499), .Z(pipeline_md_result_muxed[13]) );
  MUX2_X2 U13340 ( .A(pipeline_md_resp_result[12]), .B(pipeline_md_a[12]), .S(
        n9500), .Z(pipeline_md_result_muxed[12]) );
  MUX2_X2 U13341 ( .A(pipeline_md_resp_result[11]), .B(pipeline_md_a[11]), .S(
        n9500), .Z(pipeline_md_result_muxed[11]) );
  MUX2_X2 U13342 ( .A(pipeline_md_resp_result[10]), .B(pipeline_md_a[10]), .S(
        n9500), .Z(pipeline_md_result_muxed[10]) );
  MUX2_X2 U13343 ( .A(pipeline_md_resp_result[9]), .B(pipeline_md_a[9]), .S(
        n9500), .Z(pipeline_md_result_muxed[9]) );
  MUX2_X2 U13344 ( .A(pipeline_md_resp_result[8]), .B(pipeline_md_a[8]), .S(
        n9499), .Z(pipeline_md_result_muxed[8]) );
  MUX2_X2 U13345 ( .A(pipeline_md_resp_result[7]), .B(pipeline_md_a[7]), .S(
        n9499), .Z(pipeline_md_result_muxed[7]) );
  MUX2_X2 U13346 ( .A(pipeline_md_resp_result[6]), .B(pipeline_md_a[6]), .S(
        n9500), .Z(pipeline_md_result_muxed[6]) );
  MUX2_X2 U13347 ( .A(pipeline_md_resp_result[5]), .B(pipeline_md_a[5]), .S(
        n9500), .Z(pipeline_md_result_muxed[5]) );
  INV_X4 U13348 ( .A(pipeline_md_N255), .ZN(n12674) );
  OAI22_X2 U13349 ( .A1(n1091), .A2(n9504), .B1(n9505), .B2(n12674), .ZN(
        n12675) );
  INV_X4 U13350 ( .A(n12676), .ZN(n5656) );
  MUX2_X2 U13351 ( .A(pipeline_md_resp_result[4]), .B(pipeline_md_a[4]), .S(
        n9499), .Z(pipeline_md_result_muxed[4]) );
  MUX2_X2 U13352 ( .A(pipeline_md_resp_result[3]), .B(pipeline_md_a[3]), .S(
        n9500), .Z(pipeline_md_result_muxed[3]) );
  MUX2_X2 U13353 ( .A(pipeline_md_resp_result[2]), .B(pipeline_md_a[2]), .S(
        n9499), .Z(pipeline_md_result_muxed[2]) );
  MUX2_X2 U13354 ( .A(pipeline_md_resp_result[1]), .B(pipeline_md_a[1]), .S(
        n9499), .Z(pipeline_md_result_muxed[1]) );
  MUX2_X2 U13355 ( .A(pipeline_md_resp_result[0]), .B(pipeline_md_a[0]), .S(
        n9500), .Z(pipeline_md_result_muxed[0]) );
  INV_X4 U13356 ( .A(pipeline_md_result_muxed[62]), .ZN(n12678) );
  NOR2_X2 U13357 ( .A1(pipeline_md_N345), .A2(pipeline_md_resp_result[30]), 
        .ZN(n12677) );
  OAI22_X2 U13358 ( .A1(n12678), .A2(n6692), .B1(n12677), .B2(n6667), .ZN(
        n12679) );
  AOI221_X2 U13359 ( .B1(pipeline_md_N158), .B2(n6755), .C1(pipeline_md_N126), 
        .C2(n6754), .A(n12679), .ZN(n12682) );
  NOR2_X2 U13360 ( .A1(n13058), .A2(n6693), .ZN(n12680) );
  AOI221_X2 U13361 ( .B1(pipeline_md_N216), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[30]), .A(n12680), .ZN(n12681) );
  NAND2_X2 U13362 ( .A1(n12682), .A2(n12681), .ZN(n5623) );
  NAND2_X2 U13363 ( .A1(n7183), .A2(n9521), .ZN(n13031) );
  INV_X4 U13364 ( .A(n13031), .ZN(n13034) );
  NAND2_X2 U13365 ( .A1(n13034), .A2(n12683), .ZN(n12687) );
  INV_X4 U13366 ( .A(n12683), .ZN(n12684) );
  NAND2_X2 U13367 ( .A1(pipeline_md_N94), .A2(n6797), .ZN(n12685) );
  OAI221_X2 U13368 ( .B1(n12686), .B2(n12687), .C1(n1085), .C2(n9521), .A(
        n12685), .ZN(n5718) );
  OAI22_X2 U13369 ( .A1(n1085), .A2(n9518), .B1(n1084), .B2(n9520), .ZN(n12688) );
  AOI221_X2 U13370 ( .B1(pipeline_md_N93), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[30]), .A(n12688), .ZN(n12689) );
  INV_X4 U13371 ( .A(n12689), .ZN(n5719) );
  OAI22_X2 U13372 ( .A1(n1084), .A2(n9518), .B1(n1083), .B2(n9521), .ZN(n12690) );
  AOI221_X2 U13373 ( .B1(pipeline_md_N92), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[29]), .A(n12690), .ZN(n12691) );
  INV_X4 U13374 ( .A(n12691), .ZN(n5720) );
  OAI22_X2 U13375 ( .A1(n1083), .A2(n9518), .B1(n1082), .B2(n9520), .ZN(n12692) );
  AOI221_X2 U13376 ( .B1(pipeline_md_N91), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[28]), .A(n12692), .ZN(n12693) );
  INV_X4 U13377 ( .A(n12693), .ZN(n5721) );
  OAI22_X2 U13378 ( .A1(n1082), .A2(n9518), .B1(n1081), .B2(n9521), .ZN(n12694) );
  AOI221_X2 U13379 ( .B1(pipeline_md_N90), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[27]), .A(n12694), .ZN(n12695) );
  INV_X4 U13380 ( .A(n12695), .ZN(n5722) );
  OAI22_X2 U13381 ( .A1(n1081), .A2(n9518), .B1(n1080), .B2(n9520), .ZN(n12696) );
  AOI221_X2 U13382 ( .B1(pipeline_md_N89), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[26]), .A(n12696), .ZN(n12697) );
  INV_X4 U13383 ( .A(n12697), .ZN(n5723) );
  OAI22_X2 U13384 ( .A1(n1080), .A2(n9518), .B1(n1079), .B2(n9521), .ZN(n12698) );
  AOI221_X2 U13385 ( .B1(pipeline_md_N88), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[25]), .A(n12698), .ZN(n12699) );
  INV_X4 U13386 ( .A(n12699), .ZN(n5724) );
  OAI22_X2 U13387 ( .A1(n1079), .A2(n9518), .B1(n1078), .B2(n9520), .ZN(n12700) );
  AOI221_X2 U13388 ( .B1(pipeline_md_N87), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[24]), .A(n12700), .ZN(n12701) );
  INV_X4 U13389 ( .A(n12701), .ZN(n5725) );
  OAI22_X2 U13390 ( .A1(n1078), .A2(n9518), .B1(n1077), .B2(n9521), .ZN(n12702) );
  AOI221_X2 U13391 ( .B1(pipeline_md_N86), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[23]), .A(n12702), .ZN(n12703) );
  INV_X4 U13392 ( .A(n12703), .ZN(n5726) );
  OAI22_X2 U13393 ( .A1(n1077), .A2(n9518), .B1(n1076), .B2(n9520), .ZN(n12704) );
  AOI221_X2 U13394 ( .B1(pipeline_md_N85), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[22]), .A(n12704), .ZN(n12705) );
  INV_X4 U13395 ( .A(n12705), .ZN(n5727) );
  OAI22_X2 U13396 ( .A1(n1076), .A2(n9518), .B1(n1075), .B2(n9521), .ZN(n12706) );
  AOI221_X2 U13397 ( .B1(pipeline_md_N84), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[21]), .A(n12706), .ZN(n12707) );
  INV_X4 U13398 ( .A(n12707), .ZN(n5728) );
  OAI22_X2 U13399 ( .A1(n1075), .A2(n9518), .B1(n1074), .B2(n9520), .ZN(n12708) );
  AOI221_X2 U13400 ( .B1(pipeline_md_N83), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[20]), .A(n12708), .ZN(n12709) );
  INV_X4 U13401 ( .A(n12709), .ZN(n5729) );
  OAI22_X2 U13402 ( .A1(n1074), .A2(n9518), .B1(n1073), .B2(n9521), .ZN(n12710) );
  AOI221_X2 U13403 ( .B1(pipeline_md_N82), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[19]), .A(n12710), .ZN(n12711) );
  INV_X4 U13404 ( .A(n12711), .ZN(n5730) );
  OAI22_X2 U13405 ( .A1(n1073), .A2(n9518), .B1(n1072), .B2(n9520), .ZN(n12712) );
  AOI221_X2 U13406 ( .B1(pipeline_md_N81), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[18]), .A(n12712), .ZN(n12713) );
  INV_X4 U13407 ( .A(n12713), .ZN(n5731) );
  OAI22_X2 U13408 ( .A1(n1072), .A2(n9518), .B1(n1071), .B2(n9521), .ZN(n12714) );
  AOI221_X2 U13409 ( .B1(pipeline_md_N80), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[17]), .A(n12714), .ZN(n12715) );
  INV_X4 U13410 ( .A(n12715), .ZN(n5732) );
  OAI22_X2 U13411 ( .A1(n1071), .A2(n9518), .B1(n1070), .B2(n9521), .ZN(n12716) );
  AOI221_X2 U13412 ( .B1(pipeline_md_N79), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[16]), .A(n12716), .ZN(n12717) );
  INV_X4 U13413 ( .A(n12717), .ZN(n5733) );
  OAI22_X2 U13414 ( .A1(n1070), .A2(n9518), .B1(n1069), .B2(n9520), .ZN(n12718) );
  AOI221_X2 U13415 ( .B1(pipeline_md_N78), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[15]), .A(n12718), .ZN(n12719) );
  INV_X4 U13416 ( .A(n12719), .ZN(n5734) );
  OAI22_X2 U13417 ( .A1(n1069), .A2(n13029), .B1(n1068), .B2(n9521), .ZN(
        n12720) );
  AOI221_X2 U13418 ( .B1(pipeline_md_N77), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[14]), .A(n12720), .ZN(n12721) );
  INV_X4 U13419 ( .A(n12721), .ZN(n5735) );
  OAI22_X2 U13420 ( .A1(n1068), .A2(n13029), .B1(n1067), .B2(n9520), .ZN(
        n12722) );
  AOI221_X2 U13421 ( .B1(pipeline_md_N76), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[13]), .A(n12722), .ZN(n12723) );
  INV_X4 U13422 ( .A(n12723), .ZN(n5736) );
  OAI22_X2 U13423 ( .A1(n1067), .A2(n13029), .B1(n1066), .B2(n9520), .ZN(
        n12724) );
  INV_X4 U13424 ( .A(n12725), .ZN(n5737) );
  OAI22_X2 U13425 ( .A1(n1066), .A2(n13029), .B1(n1065), .B2(n9521), .ZN(
        n12726) );
  AOI221_X2 U13426 ( .B1(pipeline_md_N74), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[11]), .A(n12726), .ZN(n12727) );
  INV_X4 U13427 ( .A(n12727), .ZN(n5738) );
  OAI22_X2 U13428 ( .A1(n1065), .A2(n13029), .B1(n1064), .B2(n9521), .ZN(
        n12728) );
  AOI221_X2 U13429 ( .B1(pipeline_md_N73), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[10]), .A(n12728), .ZN(n12729) );
  INV_X4 U13430 ( .A(n12729), .ZN(n5739) );
  OAI22_X2 U13431 ( .A1(n1064), .A2(n13029), .B1(n1063), .B2(n9521), .ZN(
        n12730) );
  AOI221_X2 U13432 ( .B1(pipeline_md_N72), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[9]), .A(n12730), .ZN(n12731) );
  INV_X4 U13433 ( .A(n12731), .ZN(n5740) );
  OAI22_X2 U13434 ( .A1(n1063), .A2(n13029), .B1(n1062), .B2(n9521), .ZN(
        n12732) );
  INV_X4 U13435 ( .A(n12733), .ZN(n5741) );
  OAI22_X2 U13436 ( .A1(n1062), .A2(n13029), .B1(n1061), .B2(n9521), .ZN(
        n12734) );
  INV_X4 U13437 ( .A(n12735), .ZN(n5742) );
  OAI22_X2 U13438 ( .A1(n1061), .A2(n9518), .B1(n1060), .B2(n9521), .ZN(n12736) );
  AOI221_X2 U13439 ( .B1(pipeline_md_N69), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[6]), .A(n12736), .ZN(n12737) );
  INV_X4 U13440 ( .A(n12737), .ZN(n5743) );
  OAI22_X2 U13441 ( .A1(n1060), .A2(n13029), .B1(n1059), .B2(n9521), .ZN(
        n12738) );
  INV_X4 U13442 ( .A(n12739), .ZN(n5744) );
  OAI22_X2 U13443 ( .A1(n1059), .A2(n13029), .B1(n1058), .B2(n9521), .ZN(
        n12740) );
  INV_X4 U13444 ( .A(n12741), .ZN(n5745) );
  OAI22_X2 U13445 ( .A1(n1058), .A2(n13029), .B1(n1057), .B2(n9521), .ZN(
        n12742) );
  INV_X4 U13446 ( .A(n12743), .ZN(n5746) );
  OAI22_X2 U13447 ( .A1(n1057), .A2(n13029), .B1(n1056), .B2(n9521), .ZN(
        n12744) );
  INV_X4 U13448 ( .A(n12745), .ZN(n5747) );
  OAI22_X2 U13449 ( .A1(n1056), .A2(n9518), .B1(n1055), .B2(n9521), .ZN(n12746) );
  INV_X4 U13450 ( .A(n12747), .ZN(n5748) );
  OAI22_X2 U13451 ( .A1(n1055), .A2(n9518), .B1(n1054), .B2(n9521), .ZN(n12748) );
  AOI221_X2 U13452 ( .B1(pipeline_md_N63), .B2(n6797), .C1(n12749), .C2(
        pipeline_rs2_data_bypassed[0]), .A(n12748), .ZN(n12750) );
  INV_X4 U13453 ( .A(n12750), .ZN(n5749) );
  OAI22_X2 U13454 ( .A1(n1053), .A2(n9521), .B1(n1054), .B2(n9518), .ZN(n5750)
         );
  OAI22_X2 U13455 ( .A1(n1052), .A2(n9520), .B1(n1053), .B2(n9518), .ZN(n5751)
         );
  OAI22_X2 U13456 ( .A1(n1051), .A2(n9521), .B1(n1052), .B2(n9518), .ZN(n5752)
         );
  OAI22_X2 U13457 ( .A1(n1050), .A2(n9520), .B1(n1051), .B2(n9518), .ZN(n5753)
         );
  OAI22_X2 U13458 ( .A1(n1049), .A2(n9521), .B1(n1050), .B2(n9518), .ZN(n5754)
         );
  OAI22_X2 U13459 ( .A1(n1048), .A2(n9520), .B1(n1049), .B2(n9518), .ZN(n5755)
         );
  OAI22_X2 U13460 ( .A1(n1047), .A2(n9521), .B1(n1048), .B2(n9518), .ZN(n5756)
         );
  OAI22_X2 U13461 ( .A1(n1046), .A2(n9520), .B1(n1047), .B2(n9518), .ZN(n5757)
         );
  OAI22_X2 U13462 ( .A1(n1045), .A2(n9521), .B1(n1046), .B2(n9518), .ZN(n5758)
         );
  OAI22_X2 U13463 ( .A1(n1044), .A2(n9520), .B1(n1045), .B2(n9518), .ZN(n5759)
         );
  OAI22_X2 U13464 ( .A1(n1043), .A2(n9520), .B1(n1044), .B2(n9518), .ZN(n5760)
         );
  OAI22_X2 U13465 ( .A1(n1042), .A2(n9520), .B1(n1043), .B2(n9518), .ZN(n5761)
         );
  OAI22_X2 U13466 ( .A1(n1041), .A2(n9520), .B1(n1042), .B2(n9518), .ZN(n5762)
         );
  OAI22_X2 U13467 ( .A1(n1040), .A2(n9520), .B1(n1041), .B2(n9518), .ZN(n5763)
         );
  OAI22_X2 U13473 ( .A1(n1034), .A2(n9520), .B1(n1035), .B2(n13029), .ZN(n5769) );
  OAI22_X2 U13474 ( .A1(n1033), .A2(n9520), .B1(n1034), .B2(n13029), .ZN(n5770) );
  OAI22_X2 U13475 ( .A1(n1032), .A2(n9520), .B1(n1033), .B2(n13029), .ZN(n5771) );
  OAI22_X2 U13476 ( .A1(n1031), .A2(n9520), .B1(n1032), .B2(n13029), .ZN(n5772) );
  OAI22_X2 U13477 ( .A1(n1030), .A2(n9521), .B1(n1031), .B2(n13029), .ZN(n5773) );
  OAI22_X2 U13478 ( .A1(n12751), .A2(n9521), .B1(n1030), .B2(n13029), .ZN(
        n5774) );
  OAI22_X2 U13479 ( .A1(n9521), .A2(n6919), .B1(n9518), .B2(n12751), .ZN(n5775) );
  OAI22_X2 U13480 ( .A1(n9521), .A2(n6718), .B1(n9518), .B2(n6919), .ZN(n5776)
         );
  OAI22_X2 U13481 ( .A1(n9521), .A2(n6760), .B1(n9518), .B2(n6718), .ZN(n5777)
         );
  OAI22_X2 U13482 ( .A1(n9521), .A2(n6920), .B1(n9518), .B2(n6760), .ZN(n5778)
         );
  OAI22_X2 U13483 ( .A1(n9521), .A2(n6759), .B1(n9518), .B2(n6920), .ZN(n5779)
         );
  OAI22_X2 U13484 ( .A1(n9521), .A2(n6921), .B1(n9518), .B2(n6759), .ZN(n5780)
         );
  INV_X4 U13485 ( .A(pipeline_md_N249), .ZN(n12752) );
  OAI22_X2 U13486 ( .A1(n9501), .A2(n12752), .B1(n960), .B2(n6809), .ZN(n5590)
         );
  INV_X4 U13487 ( .A(pipeline_md_result_muxed[63]), .ZN(n12755) );
  NOR2_X2 U13488 ( .A1(pipeline_md_N346), .A2(pipeline_md_resp_result[31]), 
        .ZN(n12754) );
  OAI22_X2 U13489 ( .A1(n12755), .A2(n6692), .B1(n12754), .B2(n6667), .ZN(
        n12756) );
  AOI221_X2 U13490 ( .B1(pipeline_md_N159), .B2(n6755), .C1(pipeline_md_N127), 
        .C2(n6754), .A(n12756), .ZN(n12759) );
  NOR2_X2 U13491 ( .A1(n13057), .A2(n6693), .ZN(n12757) );
  AOI221_X2 U13492 ( .B1(pipeline_md_N217), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[31]), .A(n12757), .ZN(n12758) );
  NAND2_X2 U13493 ( .A1(n12759), .A2(n12758), .ZN(n5622) );
  OAI22_X2 U13494 ( .A1(n7214), .A2(n6691), .B1(n470), .B2(n9525), .ZN(n6365)
         );
  INV_X4 U13495 ( .A(pipeline_md_N282), .ZN(n12760) );
  OAI22_X2 U13496 ( .A1(n13057), .A2(n9504), .B1(n9505), .B2(n12760), .ZN(
        n12761) );
  AOI221_X2 U13497 ( .B1(pipeline_md_N60), .B2(n6798), .C1(n6808), .C2(
        pipeline_rs1_data_bypassed[31]), .A(n12761), .ZN(n12762) );
  INV_X4 U13498 ( .A(n12762), .ZN(n5684) );
  INV_X4 U13499 ( .A(pipeline_md_N314), .ZN(n12764) );
  OAI22_X2 U13500 ( .A1(n9505), .A2(n12764), .B1(n1150), .B2(n9504), .ZN(n5717) );
  INV_X4 U13501 ( .A(pipeline_md_result_muxed[36]), .ZN(n12767) );
  NOR2_X2 U13502 ( .A1(pipeline_md_N319), .A2(pipeline_md_resp_result[4]), 
        .ZN(n12766) );
  OAI22_X2 U13503 ( .A1(n12767), .A2(n6692), .B1(n12766), .B2(n6667), .ZN(
        n12768) );
  AOI221_X2 U13504 ( .B1(pipeline_md_N132), .B2(n6755), .C1(pipeline_md_N100), 
        .C2(n6754), .A(n12768), .ZN(n12771) );
  NOR2_X2 U13505 ( .A1(n1091), .A2(n6693), .ZN(n12769) );
  AOI221_X2 U13506 ( .B1(pipeline_md_N190), .B2(n9502), .C1(n6699), .C2(
        pipeline_md_resp_result[4]), .A(n12769), .ZN(n12770) );
  NAND2_X2 U13507 ( .A1(n12771), .A2(n12770), .ZN(n5649) );
  INV_X4 U13508 ( .A(n12772), .ZN(n12790) );
  INV_X4 U13509 ( .A(n12773), .ZN(n12781) );
  OAI22_X2 U13510 ( .A1(n12777), .A2(n12776), .B1(n12775), .B2(n12774), .ZN(
        n12778) );
  AOI221_X2 U13511 ( .B1(n9511), .B2(n12781), .C1(n12780), .C2(n12779), .A(
        n12778), .ZN(n12782) );
  INV_X4 U13512 ( .A(n12782), .ZN(n12789) );
  NAND2_X2 U13513 ( .A1(n9479), .A2(n12800), .ZN(n12784) );
  NAND2_X2 U13514 ( .A1(n12784), .A2(n12783), .ZN(n12788) );
  NOR2_X2 U13515 ( .A1(n6803), .A2(n12791), .ZN(n12798) );
  MUX2_X2 U13516 ( .A(n12793), .B(n9479), .S(n12792), .Z(n12797) );
  NOR2_X2 U13517 ( .A1(n12795), .A2(n12794), .ZN(n12796) );
  NOR4_X2 U13518 ( .A1(n12798), .A2(n12797), .A3(n9513), .A4(n12796), .ZN(
        n12799) );
  NOR2_X2 U13519 ( .A1(n12800), .A2(n12799), .ZN(n12801) );
  AOI221_X2 U13520 ( .B1(pipeline_alu_N257), .B2(n6812), .C1(pipeline_alu_N63), 
        .C2(n6813), .A(n12801), .ZN(n12802) );
  NAND2_X2 U13521 ( .A1(n12803), .A2(n12802), .ZN(dmem_haddr[4]) );
  MUX2_X2 U13522 ( .A(pipeline_alu_out_WB[4]), .B(dmem_haddr[4]), .S(n9523), 
        .Z(n5840) );
  OAI22_X2 U13523 ( .A1(n1905), .A2(n12806), .B1(n9515), .B2(n12804), .ZN(
        n12807) );
  AOI221_X2 U13524 ( .B1(pipeline_alu_out_WB[4]), .B2(n12809), .C1(n6670), 
        .C2(n12808), .A(n12807), .ZN(n12810) );
  INV_X4 U13525 ( .A(n12810), .ZN(n5808) );
  OAI22_X2 U13526 ( .A1(n1519), .A2(n6660), .B1(n1905), .B2(n9516), .ZN(n6211)
         );
  OAI22_X2 U13527 ( .A1(n6713), .A2(n6691), .B1(n416), .B2(n9524), .ZN(n6338)
         );
  NAND2_X2 U13528 ( .A1(n12811), .A2(pipeline_ctrl_N81), .ZN(n12812) );
  OAI221_X2 U13529 ( .B1(n12815), .B2(n12816), .C1(n1905), .C2(n12820), .A(
        n12812), .ZN(n5981) );
  NOR2_X2 U13530 ( .A1(n10323), .A2(n12816), .ZN(n12813) );
  NOR2_X2 U13531 ( .A1(n12813), .A2(n12817), .ZN(n12814) );
  OAI221_X2 U13532 ( .B1(n12815), .B2(n12822), .C1(n1911), .C2(n12820), .A(
        n12814), .ZN(n6298) );
  NOR2_X2 U13533 ( .A1(n10407), .A2(n12816), .ZN(n12818) );
  NOR2_X2 U13534 ( .A1(n12818), .A2(n12817), .ZN(n12819) );
  OAI221_X2 U13535 ( .B1(n12822), .B2(n12821), .C1(n1909), .C2(n12820), .A(
        n12819), .ZN(n6296) );
  INV_X4 U13536 ( .A(imem_hrdata[21]), .ZN(n12824) );
  OAI22_X2 U13537 ( .A1(n12826), .A2(n12825), .B1(n9599), .B2(n12829), .ZN(
        n6207) );
  OAI22_X2 U13538 ( .A1(n787), .A2(n12829), .B1(n12828), .B2(n12827), .ZN(
        n6251) );
  AOI221_X2 U13539 ( .B1(imem_hrdata[1]), .B2(n12832), .C1(n9517), .C2(
        pipeline_inst_DX[1]), .A(n12831), .ZN(n12830) );
  INV_X4 U13540 ( .A(n12830), .ZN(n6256) );
  AOI221_X2 U13541 ( .B1(imem_hrdata[0]), .B2(n12832), .C1(n9517), .C2(
        pipeline_inst_DX[0]), .A(n12831), .ZN(n12833) );
  INV_X4 U13542 ( .A(n12833), .ZN(n6294) );
  NAND2_X2 U13543 ( .A1(n12835), .A2(n12834), .ZN(n12837) );
  NAND2_X2 U13544 ( .A1(n12837), .A2(n12836), .ZN(n12838) );
  MUX2_X2 U13545 ( .A(pipeline_wb_src_sel_WB_0_), .B(n12838), .S(n9522), .Z(
        n6255) );
  MUX2_X2 U13546 ( .A(pipeline_dmem_type_WB[2]), .B(pipeline_dmem_type_2_), 
        .S(n9524), .Z(n6276) );
  MUX2_X2 U13547 ( .A(pipeline_dmem_type_WB[1]), .B(dmem_hsize[1]), .S(n9523), 
        .Z(n6274) );
  MUX2_X2 U13548 ( .A(pipeline_dmem_type_WB[0]), .B(dmem_hsize[0]), .S(n9522), 
        .Z(n6272) );
  NAND2_X2 U13549 ( .A1(pipeline_wb_src_sel_WB_0_), .A2(n12839), .ZN(n12945)
         );
  INV_X4 U13550 ( .A(n12985), .ZN(n12898) );
  NAND2_X2 U13551 ( .A1(n12898), .A2(pipeline_dmem_type_WB[1]), .ZN(n12899) );
  NAND2_X2 U13552 ( .A1(n12896), .A2(dmem_hrdata[31]), .ZN(n12851) );
  INV_X4 U13553 ( .A(dmem_hrdata[23]), .ZN(n12869) );
  INV_X4 U13554 ( .A(dmem_hrdata[15]), .ZN(n12842) );
  INV_X4 U13555 ( .A(n12979), .ZN(n12840) );
  NAND2_X2 U13556 ( .A1(dmem_hrdata[31]), .A2(n12840), .ZN(n12841) );
  OAI221_X2 U13557 ( .B1(n12891), .B2(n12869), .C1(n9408), .C2(n12842), .A(
        n12841), .ZN(n12901) );
  NOR3_X2 U13558 ( .A1(pipeline_dmem_type_WB[1]), .A2(pipeline_dmem_type_WB[2]), .A3(n12985), .ZN(n12843) );
  NAND3_X2 U13559 ( .A1(n12901), .A2(pipeline_dmem_type_WB[0]), .A3(n12843), 
        .ZN(n12850) );
  INV_X4 U13560 ( .A(n12891), .ZN(n12984) );
  INV_X4 U13561 ( .A(dmem_hrdata[31]), .ZN(n12868) );
  OAI22_X2 U13562 ( .A1(n12981), .A2(n12868), .B1(n12979), .B2(n12869), .ZN(
        n12844) );
  AOI221_X2 U13563 ( .B1(dmem_hrdata[15]), .B2(n12984), .C1(dmem_hrdata[7]), 
        .C2(n12983), .A(n12844), .ZN(n12845) );
  OR2_X1 U13564 ( .A1(n12845), .A2(n12985), .ZN(n12946) );
  INV_X4 U13565 ( .A(n12946), .ZN(n12849) );
  INV_X4 U13566 ( .A(n12893), .ZN(n12865) );
  MUX2_X2 U13567 ( .A(pipeline_regfile_data[1023]), .B(n9412), .S(n6673), .Z(
        n4628) );
  NAND2_X2 U13568 ( .A1(n12896), .A2(dmem_hrdata[30]), .ZN(n12853) );
  MUX2_X2 U13569 ( .A(pipeline_regfile_data[1022]), .B(n9413), .S(n6673), .Z(
        n4659) );
  NAND2_X2 U13570 ( .A1(n12896), .A2(dmem_hrdata[29]), .ZN(n12855) );
  MUX2_X2 U13571 ( .A(pipeline_regfile_data[1021]), .B(n9414), .S(n6673), .Z(
        n4690) );
  NAND2_X2 U13572 ( .A1(n12896), .A2(dmem_hrdata[28]), .ZN(n12857) );
  MUX2_X2 U13573 ( .A(pipeline_regfile_data[1020]), .B(n9415), .S(n6673), .Z(
        n4721) );
  NAND2_X2 U13574 ( .A1(n12896), .A2(dmem_hrdata[27]), .ZN(n12859) );
  MUX2_X2 U13575 ( .A(pipeline_regfile_data[1019]), .B(n9416), .S(n6673), .Z(
        n4752) );
  NAND2_X2 U13576 ( .A1(n12896), .A2(dmem_hrdata[26]), .ZN(n12861) );
  MUX2_X2 U13577 ( .A(pipeline_regfile_data[1018]), .B(n9417), .S(n6673), .Z(
        n4783) );
  NAND2_X2 U13578 ( .A1(n12896), .A2(dmem_hrdata[25]), .ZN(n12863) );
  MUX2_X2 U13579 ( .A(pipeline_regfile_data[1017]), .B(n9418), .S(n6673), .Z(
        n4814) );
  NAND2_X2 U13580 ( .A1(n12896), .A2(dmem_hrdata[24]), .ZN(n12866) );
  MUX2_X2 U13581 ( .A(pipeline_regfile_data[1016]), .B(n9419), .S(n6673), .Z(
        n4845) );
  OAI22_X2 U13582 ( .A1(n9408), .A2(n12869), .B1(n12891), .B2(n12868), .ZN(
        n12871) );
  AOI221_X2 U13583 ( .B1(n12896), .B2(n12871), .C1(n12945), .C2(n12870), .A(
        n12893), .ZN(n12872) );
  INV_X4 U13584 ( .A(n12872), .ZN(n13005) );
  MUX2_X2 U13585 ( .A(pipeline_regfile_data[1015]), .B(n13005), .S(n6673), .Z(
        n4876) );
  INV_X4 U13586 ( .A(dmem_hrdata[22]), .ZN(n12948) );
  INV_X4 U13587 ( .A(dmem_hrdata[30]), .ZN(n12949) );
  OAI22_X2 U13588 ( .A1(n9408), .A2(n12948), .B1(n12891), .B2(n12949), .ZN(
        n12874) );
  AOI221_X2 U13589 ( .B1(n12896), .B2(n12874), .C1(n12945), .C2(n12873), .A(
        n12893), .ZN(n12875) );
  INV_X4 U13590 ( .A(n12875), .ZN(n13006) );
  MUX2_X2 U13591 ( .A(pipeline_regfile_data[1014]), .B(n13006), .S(n6673), .Z(
        n4907) );
  INV_X4 U13592 ( .A(dmem_hrdata[21]), .ZN(n12953) );
  INV_X4 U13593 ( .A(dmem_hrdata[29]), .ZN(n12954) );
  OAI22_X2 U13594 ( .A1(n9408), .A2(n12953), .B1(n12891), .B2(n12954), .ZN(
        n12877) );
  AOI221_X2 U13595 ( .B1(n12896), .B2(n12877), .C1(n12945), .C2(n12876), .A(
        n12893), .ZN(n12878) );
  INV_X4 U13596 ( .A(n12878), .ZN(n13007) );
  MUX2_X2 U13597 ( .A(pipeline_regfile_data[1013]), .B(n13007), .S(n6673), .Z(
        n4938) );
  INV_X4 U13598 ( .A(dmem_hrdata[20]), .ZN(n12958) );
  INV_X4 U13599 ( .A(dmem_hrdata[28]), .ZN(n12959) );
  OAI22_X2 U13600 ( .A1(n9409), .A2(n12958), .B1(n12891), .B2(n12959), .ZN(
        n12880) );
  AOI221_X2 U13601 ( .B1(n12896), .B2(n12880), .C1(n12945), .C2(n12879), .A(
        n12893), .ZN(n12881) );
  INV_X4 U13602 ( .A(n12881), .ZN(n13008) );
  MUX2_X2 U13603 ( .A(pipeline_regfile_data[1012]), .B(n13008), .S(n6673), .Z(
        n4969) );
  INV_X4 U13604 ( .A(dmem_hrdata[19]), .ZN(n12963) );
  INV_X4 U13605 ( .A(dmem_hrdata[27]), .ZN(n12964) );
  OAI22_X2 U13606 ( .A1(n9408), .A2(n12963), .B1(n12891), .B2(n12964), .ZN(
        n12883) );
  AOI221_X2 U13607 ( .B1(n12896), .B2(n12883), .C1(n12945), .C2(n12882), .A(
        n12893), .ZN(n12884) );
  INV_X4 U13608 ( .A(n12884), .ZN(n13009) );
  MUX2_X2 U13609 ( .A(pipeline_regfile_data[1011]), .B(n13009), .S(n6673), .Z(
        n5000) );
  INV_X4 U13610 ( .A(dmem_hrdata[18]), .ZN(n12968) );
  INV_X4 U13611 ( .A(dmem_hrdata[26]), .ZN(n12969) );
  OAI22_X2 U13612 ( .A1(n9409), .A2(n12968), .B1(n12891), .B2(n12969), .ZN(
        n12886) );
  AOI221_X2 U13613 ( .B1(n12896), .B2(n12886), .C1(n12945), .C2(n12885), .A(
        n12893), .ZN(n12887) );
  INV_X4 U13614 ( .A(n12887), .ZN(n13010) );
  MUX2_X2 U13615 ( .A(pipeline_regfile_data[1010]), .B(n13010), .S(n6673), .Z(
        n5031) );
  INV_X4 U13616 ( .A(dmem_hrdata[17]), .ZN(n12973) );
  INV_X4 U13617 ( .A(dmem_hrdata[25]), .ZN(n12974) );
  OAI22_X2 U13618 ( .A1(n9408), .A2(n12973), .B1(n12891), .B2(n12974), .ZN(
        n12889) );
  AOI221_X2 U13619 ( .B1(n12896), .B2(n12889), .C1(n12945), .C2(n12888), .A(
        n12893), .ZN(n12890) );
  INV_X4 U13620 ( .A(n12890), .ZN(n13011) );
  MUX2_X2 U13621 ( .A(pipeline_regfile_data[1009]), .B(n13011), .S(n6673), .Z(
        n5062) );
  INV_X4 U13622 ( .A(dmem_hrdata[16]), .ZN(n12978) );
  INV_X4 U13623 ( .A(dmem_hrdata[24]), .ZN(n12980) );
  OAI22_X2 U13624 ( .A1(n12978), .A2(n9409), .B1(n12980), .B2(n12891), .ZN(
        n12895) );
  AOI221_X2 U13625 ( .B1(n12896), .B2(n12895), .C1(n12945), .C2(n12894), .A(
        n12893), .ZN(n12897) );
  INV_X4 U13626 ( .A(n12897), .ZN(n13012) );
  MUX2_X2 U13627 ( .A(pipeline_regfile_data[1008]), .B(n13012), .S(n6673), .Z(
        n5093) );
  NAND2_X2 U13628 ( .A1(n12898), .A2(pipeline_dmem_type_WB[0]), .ZN(n12900) );
  NAND2_X2 U13629 ( .A1(n12900), .A2(n12899), .ZN(n12905) );
  INV_X4 U13630 ( .A(n12905), .ZN(n12903) );
  INV_X4 U13631 ( .A(n12901), .ZN(n12902) );
  MUX2_X2 U13632 ( .A(pipeline_regfile_data[1007]), .B(n9420), .S(n6673), .Z(
        n5124) );
  OAI22_X2 U13633 ( .A1(dmem_hrdata[22]), .A2(n12937), .B1(dmem_hrdata[30]), 
        .B2(n12936), .ZN(n12910) );
  INV_X4 U13634 ( .A(dmem_hrdata[14]), .ZN(n12906) );
  NAND2_X2 U13635 ( .A1(n12983), .A2(n12906), .ZN(n12907) );
  NAND2_X2 U13636 ( .A1(n6848), .A2(n12907), .ZN(n12909) );
  MUX2_X2 U13637 ( .A(pipeline_regfile_data[1006]), .B(n9421), .S(n6673), .Z(
        n5155) );
  OAI22_X2 U13638 ( .A1(dmem_hrdata[21]), .A2(n12937), .B1(dmem_hrdata[29]), 
        .B2(n12936), .ZN(n12915) );
  INV_X4 U13639 ( .A(dmem_hrdata[13]), .ZN(n12911) );
  NAND2_X2 U13640 ( .A1(n12983), .A2(n12911), .ZN(n12912) );
  NAND2_X2 U13641 ( .A1(n6848), .A2(n12912), .ZN(n12914) );
  MUX2_X2 U13642 ( .A(pipeline_regfile_data[1005]), .B(n9422), .S(n6673), .Z(
        n5186) );
  OAI22_X2 U13643 ( .A1(dmem_hrdata[20]), .A2(n12937), .B1(dmem_hrdata[28]), 
        .B2(n12936), .ZN(n12920) );
  INV_X4 U13644 ( .A(dmem_hrdata[12]), .ZN(n12916) );
  NAND2_X2 U13645 ( .A1(n12983), .A2(n12916), .ZN(n12917) );
  NAND2_X2 U13646 ( .A1(n6848), .A2(n12917), .ZN(n12919) );
  MUX2_X2 U13647 ( .A(pipeline_regfile_data[1004]), .B(n9423), .S(n6673), .Z(
        n5217) );
  OAI22_X2 U13648 ( .A1(dmem_hrdata[19]), .A2(n12937), .B1(dmem_hrdata[27]), 
        .B2(n12936), .ZN(n12925) );
  INV_X4 U13649 ( .A(dmem_hrdata[11]), .ZN(n12921) );
  NAND2_X2 U13650 ( .A1(n12983), .A2(n12921), .ZN(n12922) );
  NAND2_X2 U13651 ( .A1(n6848), .A2(n12922), .ZN(n12924) );
  OAI221_X2 U13652 ( .B1(n12925), .B2(n12924), .C1(n12923), .C2(n9407), .A(
        n12940), .ZN(n13017) );
  MUX2_X2 U13653 ( .A(pipeline_regfile_data[1003]), .B(n9424), .S(n6673), .Z(
        n5248) );
  OAI22_X2 U13654 ( .A1(dmem_hrdata[18]), .A2(n12937), .B1(dmem_hrdata[26]), 
        .B2(n12936), .ZN(n12930) );
  INV_X4 U13655 ( .A(dmem_hrdata[10]), .ZN(n12926) );
  NAND2_X2 U13656 ( .A1(n12983), .A2(n12926), .ZN(n12927) );
  NAND2_X2 U13657 ( .A1(n6848), .A2(n12927), .ZN(n12929) );
  OAI221_X2 U13658 ( .B1(n12930), .B2(n12929), .C1(n12928), .C2(n9407), .A(
        n9410), .ZN(n13018) );
  MUX2_X2 U13659 ( .A(pipeline_regfile_data[1002]), .B(n9426), .S(n6673), .Z(
        n5279) );
  OAI22_X2 U13660 ( .A1(dmem_hrdata[17]), .A2(n12937), .B1(dmem_hrdata[25]), 
        .B2(n12936), .ZN(n12935) );
  INV_X4 U13661 ( .A(dmem_hrdata[9]), .ZN(n12931) );
  NAND2_X2 U13662 ( .A1(n12983), .A2(n12931), .ZN(n12932) );
  NAND2_X2 U13663 ( .A1(n6848), .A2(n12932), .ZN(n12934) );
  OAI221_X2 U13664 ( .B1(n12935), .B2(n12934), .C1(n12933), .C2(n9407), .A(
        n9411), .ZN(n13019) );
  MUX2_X2 U13665 ( .A(pipeline_regfile_data[1001]), .B(n9428), .S(n6673), .Z(
        n5310) );
  OAI22_X2 U13666 ( .A1(dmem_hrdata[16]), .A2(n12937), .B1(dmem_hrdata[24]), 
        .B2(n12936), .ZN(n12943) );
  INV_X4 U13667 ( .A(dmem_hrdata[8]), .ZN(n12938) );
  NAND2_X2 U13668 ( .A1(n12983), .A2(n12938), .ZN(n12939) );
  NAND2_X2 U13669 ( .A1(n6848), .A2(n12939), .ZN(n12942) );
  OAI221_X2 U13670 ( .B1(n12943), .B2(n12942), .C1(n12941), .C2(n9407), .A(
        n12940), .ZN(n13020) );
  MUX2_X2 U13671 ( .A(pipeline_regfile_data[1000]), .B(n9430), .S(n6673), .Z(
        n5341) );
  NAND2_X2 U13672 ( .A1(n12945), .A2(n12944), .ZN(n12947) );
  NAND2_X2 U13673 ( .A1(n12947), .A2(n12946), .ZN(n13021) );
  MUX2_X2 U13674 ( .A(pipeline_regfile_data[999]), .B(n13021), .S(n6673), .Z(
        n5372) );
  OAI22_X2 U13675 ( .A1(n12981), .A2(n12949), .B1(n12979), .B2(n12948), .ZN(
        n12950) );
  AOI221_X2 U13676 ( .B1(dmem_hrdata[14]), .B2(n12984), .C1(dmem_hrdata[6]), 
        .C2(n12983), .A(n12950), .ZN(n12951) );
  OAI22_X2 U13677 ( .A1(n12952), .A2(n9407), .B1(n12951), .B2(n12985), .ZN(
        n13022) );
  MUX2_X2 U13678 ( .A(pipeline_regfile_data[998]), .B(n9432), .S(n6673), .Z(
        n5403) );
  OAI22_X2 U13679 ( .A1(n12981), .A2(n12954), .B1(n12979), .B2(n12953), .ZN(
        n12955) );
  AOI221_X2 U13680 ( .B1(dmem_hrdata[13]), .B2(n12984), .C1(dmem_hrdata[5]), 
        .C2(n12983), .A(n12955), .ZN(n12956) );
  OAI22_X2 U13681 ( .A1(n12957), .A2(n9407), .B1(n12956), .B2(n12985), .ZN(
        n13023) );
  MUX2_X2 U13682 ( .A(pipeline_regfile_data[997]), .B(n9433), .S(n6673), .Z(
        n5434) );
  OAI22_X2 U13683 ( .A1(n12981), .A2(n12959), .B1(n12979), .B2(n12958), .ZN(
        n12960) );
  AOI221_X2 U13684 ( .B1(dmem_hrdata[12]), .B2(n12984), .C1(dmem_hrdata[4]), 
        .C2(n12983), .A(n12960), .ZN(n12961) );
  OAI22_X2 U13685 ( .A1(n12962), .A2(n9407), .B1(n12961), .B2(n12985), .ZN(
        n13024) );
  MUX2_X2 U13686 ( .A(pipeline_regfile_data[996]), .B(n9434), .S(n6673), .Z(
        n5465) );
  OAI22_X2 U13687 ( .A1(n12981), .A2(n12964), .B1(n12979), .B2(n12963), .ZN(
        n12965) );
  AOI221_X2 U13688 ( .B1(dmem_hrdata[11]), .B2(n12984), .C1(dmem_hrdata[3]), 
        .C2(n12983), .A(n12965), .ZN(n12966) );
  OAI22_X2 U13689 ( .A1(n12967), .A2(n9407), .B1(n12966), .B2(n12985), .ZN(
        n13025) );
  MUX2_X2 U13690 ( .A(pipeline_regfile_data[995]), .B(n9435), .S(n6673), .Z(
        n5496) );
  OAI22_X2 U13691 ( .A1(n12981), .A2(n12969), .B1(n12979), .B2(n12968), .ZN(
        n12970) );
  AOI221_X2 U13692 ( .B1(dmem_hrdata[10]), .B2(n12984), .C1(dmem_hrdata[2]), 
        .C2(n12983), .A(n12970), .ZN(n12971) );
  OAI22_X2 U13693 ( .A1(n12972), .A2(n9407), .B1(n12971), .B2(n12985), .ZN(
        n13026) );
  MUX2_X2 U13694 ( .A(pipeline_regfile_data[994]), .B(n9436), .S(n6673), .Z(
        n5527) );
  OAI22_X2 U13695 ( .A1(n12981), .A2(n12974), .B1(n12979), .B2(n12973), .ZN(
        n12975) );
  AOI221_X2 U13696 ( .B1(dmem_hrdata[9]), .B2(n12984), .C1(dmem_hrdata[1]), 
        .C2(n12983), .A(n12975), .ZN(n12976) );
  OAI22_X2 U13697 ( .A1(n12977), .A2(n9407), .B1(n12976), .B2(n12985), .ZN(
        n13027) );
  MUX2_X2 U13698 ( .A(pipeline_regfile_data[993]), .B(n9437), .S(n6673), .Z(
        n5558) );
  OAI22_X2 U13699 ( .A1(n12981), .A2(n12980), .B1(n12979), .B2(n12978), .ZN(
        n12982) );
  AOI221_X2 U13700 ( .B1(dmem_hrdata[8]), .B2(n12984), .C1(dmem_hrdata[0]), 
        .C2(n12983), .A(n12982), .ZN(n12986) );
  OAI22_X2 U13701 ( .A1(n12987), .A2(n9407), .B1(n12986), .B2(n12985), .ZN(
        n13028) );
  MUX2_X2 U13702 ( .A(pipeline_regfile_data[992]), .B(n9438), .S(n6673), .Z(
        n5589) );
  MUX2_X2 U13703 ( .A(pipeline_regfile_data[991]), .B(n12997), .S(n6674), .Z(
        n4627) );
  MUX2_X2 U13704 ( .A(pipeline_regfile_data[990]), .B(n12998), .S(n6674), .Z(
        n4658) );
  MUX2_X2 U13705 ( .A(pipeline_regfile_data[989]), .B(n12999), .S(n6674), .Z(
        n4689) );
  MUX2_X2 U13706 ( .A(pipeline_regfile_data[988]), .B(n13000), .S(n6674), .Z(
        n4720) );
  MUX2_X2 U13707 ( .A(pipeline_regfile_data[987]), .B(n13001), .S(n6674), .Z(
        n4751) );
  MUX2_X2 U13708 ( .A(pipeline_regfile_data[986]), .B(n13002), .S(n6674), .Z(
        n4782) );
  MUX2_X2 U13709 ( .A(pipeline_regfile_data[985]), .B(n13003), .S(n6674), .Z(
        n4813) );
  MUX2_X2 U13710 ( .A(pipeline_regfile_data[984]), .B(n13004), .S(n6674), .Z(
        n4844) );
  MUX2_X2 U13711 ( .A(pipeline_regfile_data[983]), .B(n13005), .S(n6674), .Z(
        n4875) );
  MUX2_X2 U13712 ( .A(pipeline_regfile_data[982]), .B(n13006), .S(n6674), .Z(
        n4906) );
  MUX2_X2 U13713 ( .A(pipeline_regfile_data[981]), .B(n13007), .S(n6674), .Z(
        n4937) );
  MUX2_X2 U13714 ( .A(pipeline_regfile_data[980]), .B(n13008), .S(n6674), .Z(
        n4968) );
  MUX2_X2 U13715 ( .A(pipeline_regfile_data[979]), .B(n13009), .S(n6674), .Z(
        n4999) );
  MUX2_X2 U13716 ( .A(pipeline_regfile_data[978]), .B(n13010), .S(n6674), .Z(
        n5030) );
  MUX2_X2 U13717 ( .A(pipeline_regfile_data[977]), .B(n13011), .S(n6674), .Z(
        n5061) );
  MUX2_X2 U13718 ( .A(pipeline_regfile_data[976]), .B(n13012), .S(n6674), .Z(
        n5092) );
  MUX2_X2 U13719 ( .A(pipeline_regfile_data[975]), .B(n13013), .S(n6674), .Z(
        n5123) );
  MUX2_X2 U13720 ( .A(pipeline_regfile_data[974]), .B(n13014), .S(n6674), .Z(
        n5154) );
  MUX2_X2 U13721 ( .A(pipeline_regfile_data[973]), .B(n13015), .S(n6674), .Z(
        n5185) );
  MUX2_X2 U13722 ( .A(pipeline_regfile_data[972]), .B(n13016), .S(n6674), .Z(
        n5216) );
  MUX2_X2 U13723 ( .A(pipeline_regfile_data[971]), .B(n9425), .S(n6674), .Z(
        n5247) );
  MUX2_X2 U13724 ( .A(pipeline_regfile_data[970]), .B(n9427), .S(n6674), .Z(
        n5278) );
  MUX2_X2 U13725 ( .A(pipeline_regfile_data[969]), .B(n9429), .S(n6674), .Z(
        n5309) );
  MUX2_X2 U13726 ( .A(pipeline_regfile_data[968]), .B(n9431), .S(n6674), .Z(
        n5340) );
  MUX2_X2 U13727 ( .A(pipeline_regfile_data[967]), .B(n13021), .S(n6674), .Z(
        n5371) );
  MUX2_X2 U13728 ( .A(pipeline_regfile_data[966]), .B(n13022), .S(n6674), .Z(
        n5402) );
  MUX2_X2 U13729 ( .A(pipeline_regfile_data[965]), .B(n13023), .S(n6674), .Z(
        n5433) );
  MUX2_X2 U13730 ( .A(pipeline_regfile_data[964]), .B(n13024), .S(n6674), .Z(
        n5464) );
  MUX2_X2 U13731 ( .A(pipeline_regfile_data[963]), .B(n13025), .S(n6674), .Z(
        n5495) );
  MUX2_X2 U13732 ( .A(pipeline_regfile_data[962]), .B(n13026), .S(n6674), .Z(
        n5526) );
  MUX2_X2 U13733 ( .A(pipeline_regfile_data[961]), .B(n13027), .S(n6674), .Z(
        n5557) );
  MUX2_X2 U13734 ( .A(pipeline_regfile_data[960]), .B(n13028), .S(n6674), .Z(
        n5588) );
  MUX2_X2 U13735 ( .A(pipeline_regfile_data[959]), .B(n9412), .S(n6675), .Z(
        n4626) );
  MUX2_X2 U13736 ( .A(pipeline_regfile_data[958]), .B(n9413), .S(n6675), .Z(
        n4657) );
  MUX2_X2 U13737 ( .A(pipeline_regfile_data[957]), .B(n9414), .S(n6675), .Z(
        n4688) );
  MUX2_X2 U13738 ( .A(pipeline_regfile_data[956]), .B(n9415), .S(n6675), .Z(
        n4719) );
  MUX2_X2 U13739 ( .A(pipeline_regfile_data[955]), .B(n9416), .S(n6675), .Z(
        n4750) );
  MUX2_X2 U13740 ( .A(pipeline_regfile_data[954]), .B(n9417), .S(n6675), .Z(
        n4781) );
  MUX2_X2 U13741 ( .A(pipeline_regfile_data[953]), .B(n9418), .S(n6675), .Z(
        n4812) );
  MUX2_X2 U13742 ( .A(pipeline_regfile_data[952]), .B(n9419), .S(n6675), .Z(
        n4843) );
  MUX2_X2 U13743 ( .A(pipeline_regfile_data[951]), .B(n13005), .S(n6675), .Z(
        n4874) );
  MUX2_X2 U13744 ( .A(pipeline_regfile_data[950]), .B(n13006), .S(n6675), .Z(
        n4905) );
  MUX2_X2 U13745 ( .A(pipeline_regfile_data[949]), .B(n13007), .S(n6675), .Z(
        n4936) );
  MUX2_X2 U13746 ( .A(pipeline_regfile_data[948]), .B(n13008), .S(n6675), .Z(
        n4967) );
  MUX2_X2 U13747 ( .A(pipeline_regfile_data[947]), .B(n13009), .S(n6675), .Z(
        n4998) );
  MUX2_X2 U13748 ( .A(pipeline_regfile_data[946]), .B(n13010), .S(n6675), .Z(
        n5029) );
  MUX2_X2 U13749 ( .A(pipeline_regfile_data[945]), .B(n13011), .S(n6675), .Z(
        n5060) );
  MUX2_X2 U13750 ( .A(pipeline_regfile_data[944]), .B(n13012), .S(n6675), .Z(
        n5091) );
  MUX2_X2 U13751 ( .A(pipeline_regfile_data[943]), .B(n9420), .S(n6675), .Z(
        n5122) );
  MUX2_X2 U13752 ( .A(pipeline_regfile_data[942]), .B(n9421), .S(n6675), .Z(
        n5153) );
  MUX2_X2 U13753 ( .A(pipeline_regfile_data[941]), .B(n9422), .S(n6675), .Z(
        n5184) );
  MUX2_X2 U13754 ( .A(pipeline_regfile_data[940]), .B(n9423), .S(n6675), .Z(
        n5215) );
  MUX2_X2 U13755 ( .A(pipeline_regfile_data[939]), .B(n13017), .S(n6675), .Z(
        n5246) );
  MUX2_X2 U13756 ( .A(pipeline_regfile_data[938]), .B(n13018), .S(n6675), .Z(
        n5277) );
  MUX2_X2 U13757 ( .A(pipeline_regfile_data[937]), .B(n13019), .S(n6675), .Z(
        n5308) );
  MUX2_X2 U13758 ( .A(pipeline_regfile_data[936]), .B(n13020), .S(n6675), .Z(
        n5339) );
  MUX2_X2 U13759 ( .A(pipeline_regfile_data[935]), .B(n13021), .S(n6675), .Z(
        n5370) );
  MUX2_X2 U13760 ( .A(pipeline_regfile_data[934]), .B(n9432), .S(n6675), .Z(
        n5401) );
  MUX2_X2 U13761 ( .A(pipeline_regfile_data[933]), .B(n9433), .S(n6675), .Z(
        n5432) );
  MUX2_X2 U13762 ( .A(pipeline_regfile_data[932]), .B(n9434), .S(n6675), .Z(
        n5463) );
  MUX2_X2 U13763 ( .A(pipeline_regfile_data[931]), .B(n9435), .S(n6675), .Z(
        n5494) );
  MUX2_X2 U13764 ( .A(pipeline_regfile_data[930]), .B(n9436), .S(n6675), .Z(
        n5525) );
  MUX2_X2 U13765 ( .A(pipeline_regfile_data[929]), .B(n9437), .S(n6675), .Z(
        n5556) );
  MUX2_X2 U13766 ( .A(pipeline_regfile_data[928]), .B(n9438), .S(n6675), .Z(
        n5587) );
  MUX2_X2 U13767 ( .A(pipeline_regfile_data[927]), .B(n12997), .S(n6676), .Z(
        n4625) );
  MUX2_X2 U13768 ( .A(pipeline_regfile_data[926]), .B(n12998), .S(n6676), .Z(
        n4656) );
  MUX2_X2 U13769 ( .A(pipeline_regfile_data[925]), .B(n12999), .S(n6676), .Z(
        n4687) );
  MUX2_X2 U13770 ( .A(pipeline_regfile_data[924]), .B(n13000), .S(n6676), .Z(
        n4718) );
  MUX2_X2 U13771 ( .A(pipeline_regfile_data[923]), .B(n13001), .S(n6676), .Z(
        n4749) );
  MUX2_X2 U13772 ( .A(pipeline_regfile_data[922]), .B(n13002), .S(n6676), .Z(
        n4780) );
  MUX2_X2 U13773 ( .A(pipeline_regfile_data[921]), .B(n13003), .S(n6676), .Z(
        n4811) );
  MUX2_X2 U13774 ( .A(pipeline_regfile_data[920]), .B(n13004), .S(n6676), .Z(
        n4842) );
  MUX2_X2 U13775 ( .A(pipeline_regfile_data[919]), .B(n13005), .S(n6676), .Z(
        n4873) );
  MUX2_X2 U13776 ( .A(pipeline_regfile_data[918]), .B(n13006), .S(n6676), .Z(
        n4904) );
  MUX2_X2 U13777 ( .A(pipeline_regfile_data[917]), .B(n13007), .S(n6676), .Z(
        n4935) );
  MUX2_X2 U13778 ( .A(pipeline_regfile_data[916]), .B(n13008), .S(n6676), .Z(
        n4966) );
  MUX2_X2 U13779 ( .A(pipeline_regfile_data[915]), .B(n13009), .S(n6676), .Z(
        n4997) );
  MUX2_X2 U13780 ( .A(pipeline_regfile_data[914]), .B(n13010), .S(n6676), .Z(
        n5028) );
  MUX2_X2 U13781 ( .A(pipeline_regfile_data[913]), .B(n13011), .S(n6676), .Z(
        n5059) );
  MUX2_X2 U13782 ( .A(pipeline_regfile_data[912]), .B(n13012), .S(n6676), .Z(
        n5090) );
  MUX2_X2 U13783 ( .A(pipeline_regfile_data[911]), .B(n13013), .S(n6676), .Z(
        n5121) );
  MUX2_X2 U13784 ( .A(pipeline_regfile_data[910]), .B(n13014), .S(n6676), .Z(
        n5152) );
  MUX2_X2 U13785 ( .A(pipeline_regfile_data[909]), .B(n13015), .S(n6676), .Z(
        n5183) );
  MUX2_X2 U13786 ( .A(pipeline_regfile_data[908]), .B(n13016), .S(n6676), .Z(
        n5214) );
  MUX2_X2 U13787 ( .A(pipeline_regfile_data[907]), .B(n9424), .S(n6676), .Z(
        n5245) );
  MUX2_X2 U13788 ( .A(pipeline_regfile_data[906]), .B(n9426), .S(n6676), .Z(
        n5276) );
  MUX2_X2 U13789 ( .A(pipeline_regfile_data[905]), .B(n9428), .S(n6676), .Z(
        n5307) );
  MUX2_X2 U13790 ( .A(pipeline_regfile_data[904]), .B(n9430), .S(n6676), .Z(
        n5338) );
  MUX2_X2 U13791 ( .A(pipeline_regfile_data[903]), .B(n13021), .S(n6676), .Z(
        n5369) );
  MUX2_X2 U13792 ( .A(pipeline_regfile_data[902]), .B(n13022), .S(n6676), .Z(
        n5400) );
  MUX2_X2 U13793 ( .A(pipeline_regfile_data[901]), .B(n13023), .S(n6676), .Z(
        n5431) );
  MUX2_X2 U13794 ( .A(pipeline_regfile_data[900]), .B(n13024), .S(n6676), .Z(
        n5462) );
  MUX2_X2 U13795 ( .A(pipeline_regfile_data[899]), .B(n13025), .S(n6676), .Z(
        n5493) );
  MUX2_X2 U13796 ( .A(pipeline_regfile_data[898]), .B(n13026), .S(n6676), .Z(
        n5524) );
  MUX2_X2 U13797 ( .A(pipeline_regfile_data[897]), .B(n13027), .S(n6676), .Z(
        n5555) );
  MUX2_X2 U13798 ( .A(pipeline_regfile_data[896]), .B(n13028), .S(n6676), .Z(
        n5586) );
  MUX2_X2 U13799 ( .A(pipeline_regfile_data[895]), .B(n9412), .S(n6677), .Z(
        n4624) );
  MUX2_X2 U13800 ( .A(pipeline_regfile_data[894]), .B(n9413), .S(n6677), .Z(
        n4655) );
  MUX2_X2 U13801 ( .A(pipeline_regfile_data[893]), .B(n9414), .S(n6677), .Z(
        n4686) );
  MUX2_X2 U13802 ( .A(pipeline_regfile_data[892]), .B(n9415), .S(n6677), .Z(
        n4717) );
  MUX2_X2 U13803 ( .A(pipeline_regfile_data[891]), .B(n9416), .S(n6677), .Z(
        n4748) );
  MUX2_X2 U13804 ( .A(pipeline_regfile_data[890]), .B(n9417), .S(n6677), .Z(
        n4779) );
  MUX2_X2 U13805 ( .A(pipeline_regfile_data[889]), .B(n9418), .S(n6677), .Z(
        n4810) );
  MUX2_X2 U13806 ( .A(pipeline_regfile_data[888]), .B(n9419), .S(n6677), .Z(
        n4841) );
  MUX2_X2 U13807 ( .A(pipeline_regfile_data[887]), .B(n13005), .S(n6677), .Z(
        n4872) );
  MUX2_X2 U13808 ( .A(pipeline_regfile_data[886]), .B(n13006), .S(n6677), .Z(
        n4903) );
  MUX2_X2 U13809 ( .A(pipeline_regfile_data[885]), .B(n13007), .S(n6677), .Z(
        n4934) );
  MUX2_X2 U13810 ( .A(pipeline_regfile_data[884]), .B(n13008), .S(n6677), .Z(
        n4965) );
  MUX2_X2 U13811 ( .A(pipeline_regfile_data[883]), .B(n13009), .S(n6677), .Z(
        n4996) );
  MUX2_X2 U13812 ( .A(pipeline_regfile_data[882]), .B(n13010), .S(n6677), .Z(
        n5027) );
  MUX2_X2 U13813 ( .A(pipeline_regfile_data[881]), .B(n13011), .S(n6677), .Z(
        n5058) );
  MUX2_X2 U13814 ( .A(pipeline_regfile_data[880]), .B(n13012), .S(n6677), .Z(
        n5089) );
  MUX2_X2 U13815 ( .A(pipeline_regfile_data[879]), .B(n9420), .S(n6677), .Z(
        n5120) );
  MUX2_X2 U13816 ( .A(pipeline_regfile_data[878]), .B(n9421), .S(n6677), .Z(
        n5151) );
  MUX2_X2 U13817 ( .A(pipeline_regfile_data[877]), .B(n9422), .S(n6677), .Z(
        n5182) );
  MUX2_X2 U13818 ( .A(pipeline_regfile_data[876]), .B(n9423), .S(n6677), .Z(
        n5213) );
  MUX2_X2 U13819 ( .A(pipeline_regfile_data[875]), .B(n9425), .S(n6677), .Z(
        n5244) );
  MUX2_X2 U13820 ( .A(pipeline_regfile_data[874]), .B(n9427), .S(n6677), .Z(
        n5275) );
  MUX2_X2 U13821 ( .A(pipeline_regfile_data[873]), .B(n9429), .S(n6677), .Z(
        n5306) );
  MUX2_X2 U13822 ( .A(pipeline_regfile_data[872]), .B(n9431), .S(n6677), .Z(
        n5337) );
  MUX2_X2 U13823 ( .A(pipeline_regfile_data[871]), .B(n13021), .S(n6677), .Z(
        n5368) );
  MUX2_X2 U13824 ( .A(pipeline_regfile_data[870]), .B(n9432), .S(n6677), .Z(
        n5399) );
  MUX2_X2 U13825 ( .A(pipeline_regfile_data[869]), .B(n9433), .S(n6677), .Z(
        n5430) );
  MUX2_X2 U13826 ( .A(pipeline_regfile_data[868]), .B(n9434), .S(n6677), .Z(
        n5461) );
  MUX2_X2 U13827 ( .A(pipeline_regfile_data[867]), .B(n9435), .S(n6677), .Z(
        n5492) );
  MUX2_X2 U13828 ( .A(pipeline_regfile_data[866]), .B(n9436), .S(n6677), .Z(
        n5523) );
  MUX2_X2 U13829 ( .A(pipeline_regfile_data[865]), .B(n9437), .S(n6677), .Z(
        n5554) );
  MUX2_X2 U13830 ( .A(pipeline_regfile_data[864]), .B(n9438), .S(n6677), .Z(
        n5585) );
  MUX2_X2 U13831 ( .A(pipeline_regfile_data[863]), .B(n12997), .S(n6678), .Z(
        n4623) );
  MUX2_X2 U13832 ( .A(pipeline_regfile_data[862]), .B(n12998), .S(n6678), .Z(
        n4654) );
  MUX2_X2 U13833 ( .A(pipeline_regfile_data[861]), .B(n12999), .S(n6678), .Z(
        n4685) );
  MUX2_X2 U13834 ( .A(pipeline_regfile_data[860]), .B(n13000), .S(n6678), .Z(
        n4716) );
  MUX2_X2 U13835 ( .A(pipeline_regfile_data[859]), .B(n13001), .S(n6678), .Z(
        n4747) );
  MUX2_X2 U13836 ( .A(pipeline_regfile_data[858]), .B(n13002), .S(n6678), .Z(
        n4778) );
  MUX2_X2 U13837 ( .A(pipeline_regfile_data[857]), .B(n13003), .S(n6678), .Z(
        n4809) );
  MUX2_X2 U13838 ( .A(pipeline_regfile_data[856]), .B(n13004), .S(n6678), .Z(
        n4840) );
  MUX2_X2 U13839 ( .A(pipeline_regfile_data[855]), .B(n13005), .S(n6678), .Z(
        n4871) );
  MUX2_X2 U13840 ( .A(pipeline_regfile_data[854]), .B(n13006), .S(n6678), .Z(
        n4902) );
  MUX2_X2 U13841 ( .A(pipeline_regfile_data[853]), .B(n13007), .S(n6678), .Z(
        n4933) );
  MUX2_X2 U13842 ( .A(pipeline_regfile_data[852]), .B(n13008), .S(n6678), .Z(
        n4964) );
  MUX2_X2 U13843 ( .A(pipeline_regfile_data[851]), .B(n13009), .S(n6678), .Z(
        n4995) );
  MUX2_X2 U13844 ( .A(pipeline_regfile_data[850]), .B(n13010), .S(n6678), .Z(
        n5026) );
  MUX2_X2 U13845 ( .A(pipeline_regfile_data[849]), .B(n13011), .S(n6678), .Z(
        n5057) );
  MUX2_X2 U13846 ( .A(pipeline_regfile_data[848]), .B(n13012), .S(n6678), .Z(
        n5088) );
  MUX2_X2 U13847 ( .A(pipeline_regfile_data[847]), .B(n13013), .S(n6678), .Z(
        n5119) );
  MUX2_X2 U13848 ( .A(pipeline_regfile_data[846]), .B(n13014), .S(n6678), .Z(
        n5150) );
  MUX2_X2 U13849 ( .A(pipeline_regfile_data[845]), .B(n13015), .S(n6678), .Z(
        n5181) );
  MUX2_X2 U13850 ( .A(pipeline_regfile_data[844]), .B(n13016), .S(n6678), .Z(
        n5212) );
  MUX2_X2 U13851 ( .A(pipeline_regfile_data[843]), .B(n13017), .S(n6678), .Z(
        n5243) );
  MUX2_X2 U13852 ( .A(pipeline_regfile_data[842]), .B(n13018), .S(n6678), .Z(
        n5274) );
  MUX2_X2 U13853 ( .A(pipeline_regfile_data[841]), .B(n13019), .S(n6678), .Z(
        n5305) );
  MUX2_X2 U13854 ( .A(pipeline_regfile_data[840]), .B(n13020), .S(n6678), .Z(
        n5336) );
  MUX2_X2 U13855 ( .A(pipeline_regfile_data[839]), .B(n13021), .S(n6678), .Z(
        n5367) );
  MUX2_X2 U13856 ( .A(pipeline_regfile_data[838]), .B(n13022), .S(n6678), .Z(
        n5398) );
  MUX2_X2 U13857 ( .A(pipeline_regfile_data[837]), .B(n13023), .S(n6678), .Z(
        n5429) );
  MUX2_X2 U13858 ( .A(pipeline_regfile_data[836]), .B(n13024), .S(n6678), .Z(
        n5460) );
  MUX2_X2 U13859 ( .A(pipeline_regfile_data[835]), .B(n13025), .S(n6678), .Z(
        n5491) );
  MUX2_X2 U13860 ( .A(pipeline_regfile_data[834]), .B(n13026), .S(n6678), .Z(
        n5522) );
  MUX2_X2 U13861 ( .A(pipeline_regfile_data[833]), .B(n13027), .S(n6678), .Z(
        n5553) );
  MUX2_X2 U13862 ( .A(pipeline_regfile_data[832]), .B(n13028), .S(n6678), .Z(
        n5584) );
  MUX2_X2 U13863 ( .A(pipeline_regfile_data[831]), .B(n9412), .S(n6679), .Z(
        n4622) );
  MUX2_X2 U13864 ( .A(pipeline_regfile_data[830]), .B(n9413), .S(n6679), .Z(
        n4653) );
  MUX2_X2 U13865 ( .A(pipeline_regfile_data[829]), .B(n9414), .S(n6679), .Z(
        n4684) );
  MUX2_X2 U13866 ( .A(pipeline_regfile_data[828]), .B(n9415), .S(n6679), .Z(
        n4715) );
  MUX2_X2 U13867 ( .A(pipeline_regfile_data[827]), .B(n9416), .S(n6679), .Z(
        n4746) );
  MUX2_X2 U13868 ( .A(pipeline_regfile_data[826]), .B(n9417), .S(n6679), .Z(
        n4777) );
  MUX2_X2 U13869 ( .A(pipeline_regfile_data[825]), .B(n9418), .S(n6679), .Z(
        n4808) );
  MUX2_X2 U13870 ( .A(pipeline_regfile_data[824]), .B(n9419), .S(n6679), .Z(
        n4839) );
  MUX2_X2 U13871 ( .A(pipeline_regfile_data[823]), .B(n13005), .S(n6679), .Z(
        n4870) );
  MUX2_X2 U13872 ( .A(pipeline_regfile_data[822]), .B(n13006), .S(n6679), .Z(
        n4901) );
  MUX2_X2 U13873 ( .A(pipeline_regfile_data[821]), .B(n13007), .S(n6679), .Z(
        n4932) );
  MUX2_X2 U13874 ( .A(pipeline_regfile_data[820]), .B(n13008), .S(n6679), .Z(
        n4963) );
  MUX2_X2 U13875 ( .A(pipeline_regfile_data[819]), .B(n13009), .S(n6679), .Z(
        n4994) );
  MUX2_X2 U13876 ( .A(pipeline_regfile_data[818]), .B(n13010), .S(n6679), .Z(
        n5025) );
  MUX2_X2 U13877 ( .A(pipeline_regfile_data[817]), .B(n13011), .S(n6679), .Z(
        n5056) );
  MUX2_X2 U13878 ( .A(pipeline_regfile_data[816]), .B(n13012), .S(n6679), .Z(
        n5087) );
  MUX2_X2 U13879 ( .A(pipeline_regfile_data[815]), .B(n9420), .S(n6679), .Z(
        n5118) );
  MUX2_X2 U13880 ( .A(pipeline_regfile_data[814]), .B(n9421), .S(n6679), .Z(
        n5149) );
  MUX2_X2 U13881 ( .A(pipeline_regfile_data[813]), .B(n9422), .S(n6679), .Z(
        n5180) );
  MUX2_X2 U13882 ( .A(pipeline_regfile_data[812]), .B(n9423), .S(n6679), .Z(
        n5211) );
  MUX2_X2 U13883 ( .A(pipeline_regfile_data[811]), .B(n9424), .S(n6679), .Z(
        n5242) );
  MUX2_X2 U13884 ( .A(pipeline_regfile_data[810]), .B(n9426), .S(n6679), .Z(
        n5273) );
  MUX2_X2 U13885 ( .A(pipeline_regfile_data[809]), .B(n9428), .S(n6679), .Z(
        n5304) );
  MUX2_X2 U13886 ( .A(pipeline_regfile_data[808]), .B(n9430), .S(n6679), .Z(
        n5335) );
  MUX2_X2 U13887 ( .A(pipeline_regfile_data[807]), .B(n13021), .S(n6679), .Z(
        n5366) );
  MUX2_X2 U13888 ( .A(pipeline_regfile_data[806]), .B(n9432), .S(n6679), .Z(
        n5397) );
  MUX2_X2 U13889 ( .A(pipeline_regfile_data[805]), .B(n9433), .S(n6679), .Z(
        n5428) );
  MUX2_X2 U13890 ( .A(pipeline_regfile_data[804]), .B(n9434), .S(n6679), .Z(
        n5459) );
  MUX2_X2 U13891 ( .A(pipeline_regfile_data[803]), .B(n9435), .S(n6679), .Z(
        n5490) );
  MUX2_X2 U13892 ( .A(pipeline_regfile_data[802]), .B(n9436), .S(n6679), .Z(
        n5521) );
  MUX2_X2 U13893 ( .A(pipeline_regfile_data[801]), .B(n9437), .S(n6679), .Z(
        n5552) );
  MUX2_X2 U13894 ( .A(pipeline_regfile_data[800]), .B(n9438), .S(n6679), .Z(
        n5583) );
  MUX2_X2 U13895 ( .A(pipeline_regfile_data[799]), .B(n12997), .S(n6680), .Z(
        n4621) );
  MUX2_X2 U13896 ( .A(pipeline_regfile_data[798]), .B(n12998), .S(n6680), .Z(
        n4652) );
  MUX2_X2 U13897 ( .A(pipeline_regfile_data[797]), .B(n12999), .S(n6680), .Z(
        n4683) );
  MUX2_X2 U13898 ( .A(pipeline_regfile_data[796]), .B(n13000), .S(n6680), .Z(
        n4714) );
  MUX2_X2 U13899 ( .A(pipeline_regfile_data[795]), .B(n13001), .S(n6680), .Z(
        n4745) );
  MUX2_X2 U13900 ( .A(pipeline_regfile_data[794]), .B(n13002), .S(n6680), .Z(
        n4776) );
  MUX2_X2 U13901 ( .A(pipeline_regfile_data[793]), .B(n13003), .S(n6680), .Z(
        n4807) );
  MUX2_X2 U13902 ( .A(pipeline_regfile_data[792]), .B(n13004), .S(n6680), .Z(
        n4838) );
  MUX2_X2 U13903 ( .A(pipeline_regfile_data[791]), .B(n13005), .S(n6680), .Z(
        n4869) );
  MUX2_X2 U13904 ( .A(pipeline_regfile_data[790]), .B(n13006), .S(n6680), .Z(
        n4900) );
  MUX2_X2 U13905 ( .A(pipeline_regfile_data[789]), .B(n13007), .S(n6680), .Z(
        n4931) );
  MUX2_X2 U13906 ( .A(pipeline_regfile_data[788]), .B(n13008), .S(n6680), .Z(
        n4962) );
  MUX2_X2 U13907 ( .A(pipeline_regfile_data[787]), .B(n13009), .S(n6680), .Z(
        n4993) );
  MUX2_X2 U13908 ( .A(pipeline_regfile_data[786]), .B(n13010), .S(n6680), .Z(
        n5024) );
  MUX2_X2 U13909 ( .A(pipeline_regfile_data[785]), .B(n13011), .S(n6680), .Z(
        n5055) );
  MUX2_X2 U13910 ( .A(pipeline_regfile_data[784]), .B(n13012), .S(n6680), .Z(
        n5086) );
  MUX2_X2 U13911 ( .A(pipeline_regfile_data[783]), .B(n13013), .S(n6680), .Z(
        n5117) );
  MUX2_X2 U13912 ( .A(pipeline_regfile_data[782]), .B(n13014), .S(n6680), .Z(
        n5148) );
  MUX2_X2 U13913 ( .A(pipeline_regfile_data[781]), .B(n13015), .S(n6680), .Z(
        n5179) );
  MUX2_X2 U13914 ( .A(pipeline_regfile_data[780]), .B(n13016), .S(n6680), .Z(
        n5210) );
  MUX2_X2 U13915 ( .A(pipeline_regfile_data[779]), .B(n9425), .S(n6680), .Z(
        n5241) );
  MUX2_X2 U13916 ( .A(pipeline_regfile_data[778]), .B(n9427), .S(n6680), .Z(
        n5272) );
  MUX2_X2 U13917 ( .A(pipeline_regfile_data[777]), .B(n9429), .S(n6680), .Z(
        n5303) );
  MUX2_X2 U13918 ( .A(pipeline_regfile_data[776]), .B(n9431), .S(n6680), .Z(
        n5334) );
  MUX2_X2 U13919 ( .A(pipeline_regfile_data[775]), .B(n13021), .S(n6680), .Z(
        n5365) );
  MUX2_X2 U13920 ( .A(pipeline_regfile_data[774]), .B(n13022), .S(n6680), .Z(
        n5396) );
  MUX2_X2 U13921 ( .A(pipeline_regfile_data[773]), .B(n13023), .S(n6680), .Z(
        n5427) );
  MUX2_X2 U13922 ( .A(pipeline_regfile_data[772]), .B(n13024), .S(n6680), .Z(
        n5458) );
  MUX2_X2 U13923 ( .A(pipeline_regfile_data[771]), .B(n13025), .S(n6680), .Z(
        n5489) );
  MUX2_X2 U13924 ( .A(pipeline_regfile_data[770]), .B(n13026), .S(n6680), .Z(
        n5520) );
  MUX2_X2 U13925 ( .A(pipeline_regfile_data[769]), .B(n13027), .S(n6680), .Z(
        n5551) );
  MUX2_X2 U13926 ( .A(pipeline_regfile_data[768]), .B(n13028), .S(n6680), .Z(
        n5582) );
  MUX2_X2 U13927 ( .A(pipeline_regfile_data[767]), .B(n9412), .S(n6681), .Z(
        n4620) );
  MUX2_X2 U13928 ( .A(pipeline_regfile_data[766]), .B(n9413), .S(n6681), .Z(
        n4651) );
  MUX2_X2 U13929 ( .A(pipeline_regfile_data[765]), .B(n9414), .S(n6681), .Z(
        n4682) );
  MUX2_X2 U13930 ( .A(pipeline_regfile_data[764]), .B(n9415), .S(n6681), .Z(
        n4713) );
  MUX2_X2 U13931 ( .A(pipeline_regfile_data[763]), .B(n9416), .S(n6681), .Z(
        n4744) );
  MUX2_X2 U13932 ( .A(pipeline_regfile_data[762]), .B(n9417), .S(n6681), .Z(
        n4775) );
  MUX2_X2 U13933 ( .A(pipeline_regfile_data[761]), .B(n9418), .S(n6681), .Z(
        n4806) );
  MUX2_X2 U13934 ( .A(pipeline_regfile_data[760]), .B(n9419), .S(n6681), .Z(
        n4837) );
  MUX2_X2 U13935 ( .A(pipeline_regfile_data[759]), .B(n13005), .S(n6681), .Z(
        n4868) );
  MUX2_X2 U13936 ( .A(pipeline_regfile_data[758]), .B(n13006), .S(n6681), .Z(
        n4899) );
  MUX2_X2 U13937 ( .A(pipeline_regfile_data[757]), .B(n13007), .S(n6681), .Z(
        n4930) );
  MUX2_X2 U13938 ( .A(pipeline_regfile_data[756]), .B(n13008), .S(n6681), .Z(
        n4961) );
  MUX2_X2 U13939 ( .A(pipeline_regfile_data[755]), .B(n13009), .S(n6681), .Z(
        n4992) );
  MUX2_X2 U13940 ( .A(pipeline_regfile_data[754]), .B(n13010), .S(n6681), .Z(
        n5023) );
  MUX2_X2 U13941 ( .A(pipeline_regfile_data[753]), .B(n13011), .S(n6681), .Z(
        n5054) );
  MUX2_X2 U13942 ( .A(pipeline_regfile_data[752]), .B(n13012), .S(n6681), .Z(
        n5085) );
  MUX2_X2 U13943 ( .A(pipeline_regfile_data[751]), .B(n9420), .S(n6681), .Z(
        n5116) );
  MUX2_X2 U13944 ( .A(pipeline_regfile_data[750]), .B(n9421), .S(n6681), .Z(
        n5147) );
  MUX2_X2 U13945 ( .A(pipeline_regfile_data[749]), .B(n9422), .S(n6681), .Z(
        n5178) );
  MUX2_X2 U13946 ( .A(pipeline_regfile_data[748]), .B(n9423), .S(n6681), .Z(
        n5209) );
  MUX2_X2 U13947 ( .A(pipeline_regfile_data[747]), .B(n13017), .S(n6681), .Z(
        n5240) );
  MUX2_X2 U13948 ( .A(pipeline_regfile_data[746]), .B(n13018), .S(n6681), .Z(
        n5271) );
  MUX2_X2 U13949 ( .A(pipeline_regfile_data[745]), .B(n13019), .S(n6681), .Z(
        n5302) );
  MUX2_X2 U13950 ( .A(pipeline_regfile_data[744]), .B(n13020), .S(n6681), .Z(
        n5333) );
  MUX2_X2 U13951 ( .A(pipeline_regfile_data[743]), .B(n13021), .S(n6681), .Z(
        n5364) );
  MUX2_X2 U13952 ( .A(pipeline_regfile_data[742]), .B(n9432), .S(n6681), .Z(
        n5395) );
  MUX2_X2 U13953 ( .A(pipeline_regfile_data[741]), .B(n9433), .S(n6681), .Z(
        n5426) );
  MUX2_X2 U13954 ( .A(pipeline_regfile_data[740]), .B(n9434), .S(n6681), .Z(
        n5457) );
  MUX2_X2 U13955 ( .A(pipeline_regfile_data[739]), .B(n9435), .S(n6681), .Z(
        n5488) );
  MUX2_X2 U13956 ( .A(pipeline_regfile_data[738]), .B(n9436), .S(n6681), .Z(
        n5519) );
  MUX2_X2 U13957 ( .A(pipeline_regfile_data[737]), .B(n9437), .S(n6681), .Z(
        n5550) );
  MUX2_X2 U13958 ( .A(pipeline_regfile_data[736]), .B(n9438), .S(n6681), .Z(
        n5581) );
  MUX2_X2 U13959 ( .A(pipeline_regfile_data[735]), .B(n12997), .S(n6682), .Z(
        n4619) );
  MUX2_X2 U13960 ( .A(pipeline_regfile_data[734]), .B(n12998), .S(n6682), .Z(
        n4650) );
  MUX2_X2 U13961 ( .A(pipeline_regfile_data[733]), .B(n12999), .S(n6682), .Z(
        n4681) );
  MUX2_X2 U13962 ( .A(pipeline_regfile_data[732]), .B(n13000), .S(n6682), .Z(
        n4712) );
  MUX2_X2 U13963 ( .A(pipeline_regfile_data[731]), .B(n13001), .S(n6682), .Z(
        n4743) );
  MUX2_X2 U13964 ( .A(pipeline_regfile_data[730]), .B(n13002), .S(n6682), .Z(
        n4774) );
  MUX2_X2 U13965 ( .A(pipeline_regfile_data[729]), .B(n13003), .S(n6682), .Z(
        n4805) );
  MUX2_X2 U13966 ( .A(pipeline_regfile_data[728]), .B(n13004), .S(n6682), .Z(
        n4836) );
  MUX2_X2 U13967 ( .A(pipeline_regfile_data[727]), .B(n13005), .S(n6682), .Z(
        n4867) );
  MUX2_X2 U13968 ( .A(pipeline_regfile_data[726]), .B(n13006), .S(n6682), .Z(
        n4898) );
  MUX2_X2 U13969 ( .A(pipeline_regfile_data[725]), .B(n13007), .S(n6682), .Z(
        n4929) );
  MUX2_X2 U13970 ( .A(pipeline_regfile_data[724]), .B(n13008), .S(n6682), .Z(
        n4960) );
  MUX2_X2 U13971 ( .A(pipeline_regfile_data[723]), .B(n13009), .S(n6682), .Z(
        n4991) );
  MUX2_X2 U13972 ( .A(pipeline_regfile_data[722]), .B(n13010), .S(n6682), .Z(
        n5022) );
  MUX2_X2 U13973 ( .A(pipeline_regfile_data[721]), .B(n13011), .S(n6682), .Z(
        n5053) );
  MUX2_X2 U13974 ( .A(pipeline_regfile_data[720]), .B(n13012), .S(n6682), .Z(
        n5084) );
  MUX2_X2 U13975 ( .A(pipeline_regfile_data[719]), .B(n13013), .S(n6682), .Z(
        n5115) );
  MUX2_X2 U13976 ( .A(pipeline_regfile_data[718]), .B(n13014), .S(n6682), .Z(
        n5146) );
  MUX2_X2 U13977 ( .A(pipeline_regfile_data[717]), .B(n13015), .S(n6682), .Z(
        n5177) );
  MUX2_X2 U13978 ( .A(pipeline_regfile_data[716]), .B(n13016), .S(n6682), .Z(
        n5208) );
  MUX2_X2 U13979 ( .A(pipeline_regfile_data[715]), .B(n9424), .S(n6682), .Z(
        n5239) );
  MUX2_X2 U13980 ( .A(pipeline_regfile_data[714]), .B(n9426), .S(n6682), .Z(
        n5270) );
  MUX2_X2 U13981 ( .A(pipeline_regfile_data[713]), .B(n9428), .S(n6682), .Z(
        n5301) );
  MUX2_X2 U13982 ( .A(pipeline_regfile_data[712]), .B(n9430), .S(n6682), .Z(
        n5332) );
  MUX2_X2 U13983 ( .A(pipeline_regfile_data[711]), .B(n13021), .S(n6682), .Z(
        n5363) );
  MUX2_X2 U13984 ( .A(pipeline_regfile_data[710]), .B(n13022), .S(n6682), .Z(
        n5394) );
  MUX2_X2 U13985 ( .A(pipeline_regfile_data[709]), .B(n13023), .S(n6682), .Z(
        n5425) );
  MUX2_X2 U13986 ( .A(pipeline_regfile_data[708]), .B(n13024), .S(n6682), .Z(
        n5456) );
  MUX2_X2 U13987 ( .A(pipeline_regfile_data[707]), .B(n13025), .S(n6682), .Z(
        n5487) );
  MUX2_X2 U13988 ( .A(pipeline_regfile_data[706]), .B(n13026), .S(n6682), .Z(
        n5518) );
  MUX2_X2 U13989 ( .A(pipeline_regfile_data[705]), .B(n13027), .S(n6682), .Z(
        n5549) );
  MUX2_X2 U13990 ( .A(pipeline_regfile_data[704]), .B(n13028), .S(n6682), .Z(
        n5580) );
  MUX2_X2 U13991 ( .A(pipeline_regfile_data[703]), .B(n9412), .S(n6683), .Z(
        n4618) );
  MUX2_X2 U13992 ( .A(pipeline_regfile_data[702]), .B(n9413), .S(n6683), .Z(
        n4649) );
  MUX2_X2 U13993 ( .A(pipeline_regfile_data[701]), .B(n9414), .S(n6683), .Z(
        n4680) );
  MUX2_X2 U13994 ( .A(pipeline_regfile_data[700]), .B(n9415), .S(n6683), .Z(
        n4711) );
  MUX2_X2 U13995 ( .A(pipeline_regfile_data[699]), .B(n9416), .S(n6683), .Z(
        n4742) );
  MUX2_X2 U13996 ( .A(pipeline_regfile_data[698]), .B(n9417), .S(n6683), .Z(
        n4773) );
  MUX2_X2 U13997 ( .A(pipeline_regfile_data[697]), .B(n9418), .S(n6683), .Z(
        n4804) );
  MUX2_X2 U13998 ( .A(pipeline_regfile_data[696]), .B(n9419), .S(n6683), .Z(
        n4835) );
  MUX2_X2 U13999 ( .A(pipeline_regfile_data[695]), .B(n13005), .S(n6683), .Z(
        n4866) );
  MUX2_X2 U14000 ( .A(pipeline_regfile_data[694]), .B(n13006), .S(n6683), .Z(
        n4897) );
  MUX2_X2 U14001 ( .A(pipeline_regfile_data[693]), .B(n13007), .S(n6683), .Z(
        n4928) );
  MUX2_X2 U14002 ( .A(pipeline_regfile_data[692]), .B(n13008), .S(n6683), .Z(
        n4959) );
  MUX2_X2 U14003 ( .A(pipeline_regfile_data[691]), .B(n13009), .S(n6683), .Z(
        n4990) );
  MUX2_X2 U14004 ( .A(pipeline_regfile_data[690]), .B(n13010), .S(n6683), .Z(
        n5021) );
  MUX2_X2 U14005 ( .A(pipeline_regfile_data[689]), .B(n13011), .S(n6683), .Z(
        n5052) );
  MUX2_X2 U14006 ( .A(pipeline_regfile_data[688]), .B(n13012), .S(n6683), .Z(
        n5083) );
  MUX2_X2 U14007 ( .A(pipeline_regfile_data[687]), .B(n9420), .S(n6683), .Z(
        n5114) );
  MUX2_X2 U14008 ( .A(pipeline_regfile_data[686]), .B(n9421), .S(n6683), .Z(
        n5145) );
  MUX2_X2 U14009 ( .A(pipeline_regfile_data[685]), .B(n9422), .S(n6683), .Z(
        n5176) );
  MUX2_X2 U14010 ( .A(pipeline_regfile_data[684]), .B(n9423), .S(n6683), .Z(
        n5207) );
  MUX2_X2 U14011 ( .A(pipeline_regfile_data[683]), .B(n9425), .S(n6683), .Z(
        n5238) );
  MUX2_X2 U14012 ( .A(pipeline_regfile_data[682]), .B(n9427), .S(n6683), .Z(
        n5269) );
  MUX2_X2 U14013 ( .A(pipeline_regfile_data[681]), .B(n9429), .S(n6683), .Z(
        n5300) );
  MUX2_X2 U14014 ( .A(pipeline_regfile_data[680]), .B(n9431), .S(n6683), .Z(
        n5331) );
  MUX2_X2 U14015 ( .A(pipeline_regfile_data[679]), .B(n13021), .S(n6683), .Z(
        n5362) );
  MUX2_X2 U14016 ( .A(pipeline_regfile_data[678]), .B(n9432), .S(n6683), .Z(
        n5393) );
  MUX2_X2 U14017 ( .A(pipeline_regfile_data[677]), .B(n9433), .S(n6683), .Z(
        n5424) );
  MUX2_X2 U14018 ( .A(pipeline_regfile_data[676]), .B(n9434), .S(n6683), .Z(
        n5455) );
  MUX2_X2 U14019 ( .A(pipeline_regfile_data[675]), .B(n9435), .S(n6683), .Z(
        n5486) );
  MUX2_X2 U14020 ( .A(pipeline_regfile_data[674]), .B(n9436), .S(n6683), .Z(
        n5517) );
  MUX2_X2 U14021 ( .A(pipeline_regfile_data[673]), .B(n9437), .S(n6683), .Z(
        n5548) );
  MUX2_X2 U14022 ( .A(pipeline_regfile_data[672]), .B(n9438), .S(n6683), .Z(
        n5579) );
  MUX2_X2 U14023 ( .A(pipeline_regfile_data[671]), .B(n12997), .S(n6684), .Z(
        n4617) );
  MUX2_X2 U14024 ( .A(pipeline_regfile_data[670]), .B(n12998), .S(n6684), .Z(
        n4648) );
  MUX2_X2 U14025 ( .A(pipeline_regfile_data[669]), .B(n12999), .S(n6684), .Z(
        n4679) );
  MUX2_X2 U14026 ( .A(pipeline_regfile_data[668]), .B(n13000), .S(n6684), .Z(
        n4710) );
  MUX2_X2 U14027 ( .A(pipeline_regfile_data[667]), .B(n13001), .S(n6684), .Z(
        n4741) );
  MUX2_X2 U14028 ( .A(pipeline_regfile_data[666]), .B(n13002), .S(n6684), .Z(
        n4772) );
  MUX2_X2 U14029 ( .A(pipeline_regfile_data[665]), .B(n13003), .S(n6684), .Z(
        n4803) );
  MUX2_X2 U14030 ( .A(pipeline_regfile_data[664]), .B(n13004), .S(n6684), .Z(
        n4834) );
  MUX2_X2 U14031 ( .A(pipeline_regfile_data[663]), .B(n13005), .S(n6684), .Z(
        n4865) );
  MUX2_X2 U14032 ( .A(pipeline_regfile_data[662]), .B(n13006), .S(n6684), .Z(
        n4896) );
  MUX2_X2 U14033 ( .A(pipeline_regfile_data[661]), .B(n13007), .S(n6684), .Z(
        n4927) );
  MUX2_X2 U14034 ( .A(pipeline_regfile_data[660]), .B(n13008), .S(n6684), .Z(
        n4958) );
  MUX2_X2 U14035 ( .A(pipeline_regfile_data[659]), .B(n13009), .S(n6684), .Z(
        n4989) );
  MUX2_X2 U14036 ( .A(pipeline_regfile_data[658]), .B(n13010), .S(n6684), .Z(
        n5020) );
  MUX2_X2 U14037 ( .A(pipeline_regfile_data[657]), .B(n13011), .S(n6684), .Z(
        n5051) );
  MUX2_X2 U14038 ( .A(pipeline_regfile_data[656]), .B(n13012), .S(n6684), .Z(
        n5082) );
  MUX2_X2 U14039 ( .A(pipeline_regfile_data[655]), .B(n13013), .S(n6684), .Z(
        n5113) );
  MUX2_X2 U14040 ( .A(pipeline_regfile_data[654]), .B(n13014), .S(n6684), .Z(
        n5144) );
  MUX2_X2 U14041 ( .A(pipeline_regfile_data[653]), .B(n13015), .S(n6684), .Z(
        n5175) );
  MUX2_X2 U14042 ( .A(pipeline_regfile_data[652]), .B(n13016), .S(n6684), .Z(
        n5206) );
  MUX2_X2 U14043 ( .A(pipeline_regfile_data[651]), .B(n13017), .S(n6684), .Z(
        n5237) );
  MUX2_X2 U14044 ( .A(pipeline_regfile_data[650]), .B(n13018), .S(n6684), .Z(
        n5268) );
  MUX2_X2 U14045 ( .A(pipeline_regfile_data[649]), .B(n13019), .S(n6684), .Z(
        n5299) );
  MUX2_X2 U14046 ( .A(pipeline_regfile_data[648]), .B(n13020), .S(n6684), .Z(
        n5330) );
  MUX2_X2 U14047 ( .A(pipeline_regfile_data[647]), .B(n13021), .S(n6684), .Z(
        n5361) );
  MUX2_X2 U14048 ( .A(pipeline_regfile_data[646]), .B(n13022), .S(n6684), .Z(
        n5392) );
  MUX2_X2 U14049 ( .A(pipeline_regfile_data[645]), .B(n13023), .S(n6684), .Z(
        n5423) );
  MUX2_X2 U14050 ( .A(pipeline_regfile_data[644]), .B(n13024), .S(n6684), .Z(
        n5454) );
  MUX2_X2 U14051 ( .A(pipeline_regfile_data[643]), .B(n13025), .S(n6684), .Z(
        n5485) );
  MUX2_X2 U14052 ( .A(pipeline_regfile_data[642]), .B(n13026), .S(n6684), .Z(
        n5516) );
  MUX2_X2 U14053 ( .A(pipeline_regfile_data[641]), .B(n13027), .S(n6684), .Z(
        n5547) );
  MUX2_X2 U14054 ( .A(pipeline_regfile_data[640]), .B(n13028), .S(n6684), .Z(
        n5578) );
  MUX2_X2 U14055 ( .A(pipeline_regfile_data[639]), .B(n9412), .S(n6671), .Z(
        n4616) );
  MUX2_X2 U14056 ( .A(pipeline_regfile_data[638]), .B(n9413), .S(n6671), .Z(
        n4647) );
  MUX2_X2 U14057 ( .A(pipeline_regfile_data[637]), .B(n9414), .S(n6671), .Z(
        n4678) );
  MUX2_X2 U14058 ( .A(pipeline_regfile_data[636]), .B(n9415), .S(n6671), .Z(
        n4709) );
  MUX2_X2 U14059 ( .A(pipeline_regfile_data[635]), .B(n9416), .S(n6671), .Z(
        n4740) );
  MUX2_X2 U14060 ( .A(pipeline_regfile_data[634]), .B(n9417), .S(n6671), .Z(
        n4771) );
  MUX2_X2 U14061 ( .A(pipeline_regfile_data[633]), .B(n9418), .S(n6671), .Z(
        n4802) );
  MUX2_X2 U14062 ( .A(pipeline_regfile_data[632]), .B(n9419), .S(n6671), .Z(
        n4833) );
  MUX2_X2 U14063 ( .A(pipeline_regfile_data[631]), .B(n13005), .S(n6671), .Z(
        n4864) );
  MUX2_X2 U14064 ( .A(pipeline_regfile_data[630]), .B(n13006), .S(n6671), .Z(
        n4895) );
  MUX2_X2 U14065 ( .A(pipeline_regfile_data[629]), .B(n13007), .S(n6671), .Z(
        n4926) );
  MUX2_X2 U14066 ( .A(pipeline_regfile_data[628]), .B(n13008), .S(n6671), .Z(
        n4957) );
  MUX2_X2 U14067 ( .A(pipeline_regfile_data[627]), .B(n13009), .S(n6671), .Z(
        n4988) );
  MUX2_X2 U14068 ( .A(pipeline_regfile_data[626]), .B(n13010), .S(n6671), .Z(
        n5019) );
  MUX2_X2 U14069 ( .A(pipeline_regfile_data[625]), .B(n13011), .S(n6671), .Z(
        n5050) );
  MUX2_X2 U14070 ( .A(pipeline_regfile_data[624]), .B(n13012), .S(n6671), .Z(
        n5081) );
  MUX2_X2 U14071 ( .A(pipeline_regfile_data[623]), .B(n9420), .S(n6671), .Z(
        n5112) );
  MUX2_X2 U14072 ( .A(pipeline_regfile_data[622]), .B(n9421), .S(n6671), .Z(
        n5143) );
  MUX2_X2 U14073 ( .A(pipeline_regfile_data[621]), .B(n9422), .S(n6671), .Z(
        n5174) );
  MUX2_X2 U14074 ( .A(pipeline_regfile_data[619]), .B(n9424), .S(n6671), .Z(
        n5236) );
  MUX2_X2 U14075 ( .A(pipeline_regfile_data[618]), .B(n9426), .S(n6671), .Z(
        n5267) );
  MUX2_X2 U14076 ( .A(pipeline_regfile_data[617]), .B(n9428), .S(n6671), .Z(
        n5298) );
  MUX2_X2 U14077 ( .A(pipeline_regfile_data[616]), .B(n9430), .S(n6671), .Z(
        n5329) );
  MUX2_X2 U14078 ( .A(pipeline_regfile_data[615]), .B(n13021), .S(n6671), .Z(
        n5360) );
  MUX2_X2 U14079 ( .A(pipeline_regfile_data[614]), .B(n9432), .S(n6671), .Z(
        n5391) );
  MUX2_X2 U14080 ( .A(pipeline_regfile_data[613]), .B(n9433), .S(n6671), .Z(
        n5422) );
  MUX2_X2 U14081 ( .A(pipeline_regfile_data[612]), .B(n9434), .S(n6671), .Z(
        n5453) );
  MUX2_X2 U14082 ( .A(pipeline_regfile_data[611]), .B(n9435), .S(n6671), .Z(
        n5484) );
  MUX2_X2 U14083 ( .A(pipeline_regfile_data[608]), .B(n9438), .S(n6671), .Z(
        n5577) );
  MUX2_X2 U14084 ( .A(pipeline_regfile_data[607]), .B(n12997), .S(n6685), .Z(
        n4615) );
  MUX2_X2 U14085 ( .A(pipeline_regfile_data[606]), .B(n12998), .S(n6685), .Z(
        n4646) );
  MUX2_X2 U14086 ( .A(pipeline_regfile_data[605]), .B(n12999), .S(n6685), .Z(
        n4677) );
  MUX2_X2 U14087 ( .A(pipeline_regfile_data[604]), .B(n13000), .S(n6685), .Z(
        n4708) );
  MUX2_X2 U14088 ( .A(pipeline_regfile_data[603]), .B(n13001), .S(n6685), .Z(
        n4739) );
  MUX2_X2 U14089 ( .A(pipeline_regfile_data[602]), .B(n13002), .S(n6685), .Z(
        n4770) );
  MUX2_X2 U14090 ( .A(pipeline_regfile_data[601]), .B(n13003), .S(n6685), .Z(
        n4801) );
  MUX2_X2 U14091 ( .A(pipeline_regfile_data[600]), .B(n13004), .S(n6685), .Z(
        n4832) );
  MUX2_X2 U14092 ( .A(pipeline_regfile_data[599]), .B(n13005), .S(n6685), .Z(
        n4863) );
  MUX2_X2 U14093 ( .A(pipeline_regfile_data[598]), .B(n13006), .S(n6685), .Z(
        n4894) );
  MUX2_X2 U14094 ( .A(pipeline_regfile_data[597]), .B(n13007), .S(n6685), .Z(
        n4925) );
  MUX2_X2 U14095 ( .A(pipeline_regfile_data[596]), .B(n13008), .S(n6685), .Z(
        n4956) );
  MUX2_X2 U14096 ( .A(pipeline_regfile_data[595]), .B(n13009), .S(n6685), .Z(
        n4987) );
  MUX2_X2 U14097 ( .A(pipeline_regfile_data[594]), .B(n13010), .S(n6685), .Z(
        n5018) );
  MUX2_X2 U14098 ( .A(pipeline_regfile_data[593]), .B(n13011), .S(n6685), .Z(
        n5049) );
  MUX2_X2 U14099 ( .A(pipeline_regfile_data[592]), .B(n13012), .S(n6685), .Z(
        n5080) );
  MUX2_X2 U14100 ( .A(pipeline_regfile_data[591]), .B(n13013), .S(n6685), .Z(
        n5111) );
  MUX2_X2 U14101 ( .A(pipeline_regfile_data[590]), .B(n13014), .S(n6685), .Z(
        n5142) );
  MUX2_X2 U14102 ( .A(pipeline_regfile_data[589]), .B(n13015), .S(n6685), .Z(
        n5173) );
  MUX2_X2 U14103 ( .A(pipeline_regfile_data[588]), .B(n13016), .S(n6685), .Z(
        n5204) );
  MUX2_X2 U14104 ( .A(pipeline_regfile_data[587]), .B(n9425), .S(n6685), .Z(
        n5235) );
  MUX2_X2 U14105 ( .A(pipeline_regfile_data[586]), .B(n9427), .S(n6685), .Z(
        n5266) );
  MUX2_X2 U14106 ( .A(pipeline_regfile_data[585]), .B(n9429), .S(n6685), .Z(
        n5297) );
  MUX2_X2 U14107 ( .A(pipeline_regfile_data[584]), .B(n9431), .S(n6685), .Z(
        n5328) );
  MUX2_X2 U14108 ( .A(pipeline_regfile_data[583]), .B(n13021), .S(n6685), .Z(
        n5359) );
  MUX2_X2 U14109 ( .A(pipeline_regfile_data[582]), .B(n13022), .S(n6685), .Z(
        n5390) );
  MUX2_X2 U14110 ( .A(pipeline_regfile_data[581]), .B(n13023), .S(n6685), .Z(
        n5421) );
  MUX2_X2 U14111 ( .A(pipeline_regfile_data[580]), .B(n13024), .S(n6685), .Z(
        n5452) );
  MUX2_X2 U14112 ( .A(pipeline_regfile_data[579]), .B(n13025), .S(n6685), .Z(
        n5483) );
  MUX2_X2 U14113 ( .A(pipeline_regfile_data[578]), .B(n13026), .S(n6685), .Z(
        n5514) );
  MUX2_X2 U14114 ( .A(pipeline_regfile_data[577]), .B(n13027), .S(n6685), .Z(
        n5545) );
  MUX2_X2 U14115 ( .A(pipeline_regfile_data[576]), .B(n13028), .S(n6685), .Z(
        n5576) );
  MUX2_X2 U14116 ( .A(pipeline_regfile_data[575]), .B(n9412), .S(n6672), .Z(
        n4614) );
  MUX2_X2 U14117 ( .A(pipeline_regfile_data[574]), .B(n9413), .S(n6672), .Z(
        n4645) );
  MUX2_X2 U14118 ( .A(pipeline_regfile_data[573]), .B(n9414), .S(n6672), .Z(
        n4676) );
  MUX2_X2 U14119 ( .A(pipeline_regfile_data[572]), .B(n9415), .S(n6672), .Z(
        n4707) );
  MUX2_X2 U14120 ( .A(pipeline_regfile_data[571]), .B(n9416), .S(n6672), .Z(
        n4738) );
  MUX2_X2 U14121 ( .A(pipeline_regfile_data[570]), .B(n9417), .S(n6672), .Z(
        n4769) );
  MUX2_X2 U14122 ( .A(pipeline_regfile_data[569]), .B(n9418), .S(n6672), .Z(
        n4800) );
  MUX2_X2 U14123 ( .A(pipeline_regfile_data[568]), .B(n9419), .S(n6672), .Z(
        n4831) );
  MUX2_X2 U14124 ( .A(pipeline_regfile_data[567]), .B(n13005), .S(n6672), .Z(
        n4862) );
  MUX2_X2 U14125 ( .A(pipeline_regfile_data[566]), .B(n13006), .S(n6672), .Z(
        n4893) );
  MUX2_X2 U14126 ( .A(pipeline_regfile_data[565]), .B(n13007), .S(n6672), .Z(
        n4924) );
  MUX2_X2 U14127 ( .A(pipeline_regfile_data[564]), .B(n13008), .S(n6672), .Z(
        n4955) );
  MUX2_X2 U14128 ( .A(pipeline_regfile_data[563]), .B(n13009), .S(n6672), .Z(
        n4986) );
  MUX2_X2 U14129 ( .A(pipeline_regfile_data[562]), .B(n13010), .S(n6672), .Z(
        n5017) );
  MUX2_X2 U14130 ( .A(pipeline_regfile_data[561]), .B(n13011), .S(n6672), .Z(
        n5048) );
  MUX2_X2 U14131 ( .A(pipeline_regfile_data[560]), .B(n13012), .S(n6672), .Z(
        n5079) );
  MUX2_X2 U14132 ( .A(pipeline_regfile_data[559]), .B(n9420), .S(n6672), .Z(
        n5110) );
  MUX2_X2 U14133 ( .A(pipeline_regfile_data[558]), .B(n9421), .S(n6672), .Z(
        n5141) );
  MUX2_X2 U14134 ( .A(pipeline_regfile_data[557]), .B(n9422), .S(n6672), .Z(
        n5172) );
  MUX2_X2 U14135 ( .A(pipeline_regfile_data[556]), .B(n9423), .S(n6672), .Z(
        n5203) );
  MUX2_X2 U14136 ( .A(pipeline_regfile_data[555]), .B(n13017), .S(n6672), .Z(
        n5234) );
  MUX2_X2 U14137 ( .A(pipeline_regfile_data[554]), .B(n13018), .S(n6672), .Z(
        n5265) );
  MUX2_X2 U14138 ( .A(pipeline_regfile_data[553]), .B(n13019), .S(n6672), .Z(
        n5296) );
  MUX2_X2 U14139 ( .A(pipeline_regfile_data[552]), .B(n13020), .S(n6672), .Z(
        n5327) );
  MUX2_X2 U14140 ( .A(pipeline_regfile_data[551]), .B(n13021), .S(n6672), .Z(
        n5358) );
  MUX2_X2 U14141 ( .A(pipeline_regfile_data[550]), .B(n9432), .S(n6672), .Z(
        n5389) );
  MUX2_X2 U14142 ( .A(pipeline_regfile_data[549]), .B(n9433), .S(n6672), .Z(
        n5420) );
  MUX2_X2 U14143 ( .A(pipeline_regfile_data[548]), .B(n9434), .S(n6672), .Z(
        n5451) );
  MUX2_X2 U14144 ( .A(pipeline_regfile_data[547]), .B(n9435), .S(n6672), .Z(
        n5482) );
  MUX2_X2 U14145 ( .A(pipeline_regfile_data[546]), .B(n9436), .S(n6672), .Z(
        n5513) );
  MUX2_X2 U14146 ( .A(pipeline_regfile_data[544]), .B(n9438), .S(n6672), .Z(
        n5575) );
  MUX2_X2 U14147 ( .A(pipeline_regfile_data[543]), .B(n12997), .S(n6686), .Z(
        n4613) );
  MUX2_X2 U14148 ( .A(pipeline_regfile_data[542]), .B(n12998), .S(n6686), .Z(
        n4644) );
  MUX2_X2 U14149 ( .A(pipeline_regfile_data[541]), .B(n12999), .S(n6686), .Z(
        n4675) );
  MUX2_X2 U14150 ( .A(pipeline_regfile_data[540]), .B(n13000), .S(n6686), .Z(
        n4706) );
  MUX2_X2 U14151 ( .A(pipeline_regfile_data[539]), .B(n13001), .S(n6686), .Z(
        n4737) );
  MUX2_X2 U14152 ( .A(pipeline_regfile_data[538]), .B(n13002), .S(n6686), .Z(
        n4768) );
  MUX2_X2 U14153 ( .A(pipeline_regfile_data[537]), .B(n13003), .S(n6686), .Z(
        n4799) );
  MUX2_X2 U14154 ( .A(pipeline_regfile_data[536]), .B(n13004), .S(n6686), .Z(
        n4830) );
  MUX2_X2 U14155 ( .A(pipeline_regfile_data[535]), .B(n13005), .S(n6686), .Z(
        n4861) );
  MUX2_X2 U14156 ( .A(pipeline_regfile_data[534]), .B(n13006), .S(n6686), .Z(
        n4892) );
  MUX2_X2 U14157 ( .A(pipeline_regfile_data[533]), .B(n13007), .S(n6686), .Z(
        n4923) );
  MUX2_X2 U14158 ( .A(pipeline_regfile_data[532]), .B(n13008), .S(n6686), .Z(
        n4954) );
  MUX2_X2 U14159 ( .A(pipeline_regfile_data[531]), .B(n13009), .S(n6686), .Z(
        n4985) );
  MUX2_X2 U14160 ( .A(pipeline_regfile_data[530]), .B(n13010), .S(n6686), .Z(
        n5016) );
  MUX2_X2 U14161 ( .A(pipeline_regfile_data[529]), .B(n13011), .S(n6686), .Z(
        n5047) );
  MUX2_X2 U14162 ( .A(pipeline_regfile_data[528]), .B(n13012), .S(n6686), .Z(
        n5078) );
  MUX2_X2 U14163 ( .A(pipeline_regfile_data[527]), .B(n13013), .S(n6686), .Z(
        n5109) );
  MUX2_X2 U14164 ( .A(pipeline_regfile_data[526]), .B(n13014), .S(n6686), .Z(
        n5140) );
  MUX2_X2 U14165 ( .A(pipeline_regfile_data[525]), .B(n13015), .S(n6686), .Z(
        n5171) );
  MUX2_X2 U14166 ( .A(pipeline_regfile_data[524]), .B(n13016), .S(n6686), .Z(
        n5202) );
  MUX2_X2 U14167 ( .A(pipeline_regfile_data[523]), .B(n9424), .S(n6686), .Z(
        n5233) );
  MUX2_X2 U14168 ( .A(pipeline_regfile_data[522]), .B(n9426), .S(n6686), .Z(
        n5264) );
  MUX2_X2 U14169 ( .A(pipeline_regfile_data[521]), .B(n9428), .S(n6686), .Z(
        n5295) );
  MUX2_X2 U14170 ( .A(pipeline_regfile_data[520]), .B(n9430), .S(n6686), .Z(
        n5326) );
  MUX2_X2 U14171 ( .A(pipeline_regfile_data[519]), .B(n13021), .S(n6686), .Z(
        n5357) );
  MUX2_X2 U14172 ( .A(pipeline_regfile_data[518]), .B(n13022), .S(n6686), .Z(
        n5388) );
  MUX2_X2 U14173 ( .A(pipeline_regfile_data[517]), .B(n13023), .S(n6686), .Z(
        n5419) );
  MUX2_X2 U14174 ( .A(pipeline_regfile_data[516]), .B(n13024), .S(n6686), .Z(
        n5450) );
  MUX2_X2 U14175 ( .A(pipeline_regfile_data[515]), .B(n13025), .S(n6686), .Z(
        n5481) );
  MUX2_X2 U14176 ( .A(pipeline_regfile_data[514]), .B(n13026), .S(n6686), .Z(
        n5512) );
  MUX2_X2 U14177 ( .A(pipeline_regfile_data[513]), .B(n13027), .S(n6686), .Z(
        n5543) );
  MUX2_X2 U14178 ( .A(pipeline_regfile_data[512]), .B(n13028), .S(n6686), .Z(
        n5574) );
  MUX2_X2 U14179 ( .A(pipeline_regfile_data[511]), .B(n9412), .S(n6644), .Z(
        n4612) );
  MUX2_X2 U14180 ( .A(pipeline_regfile_data[510]), .B(n9413), .S(n6644), .Z(
        n4643) );
  MUX2_X2 U14181 ( .A(pipeline_regfile_data[509]), .B(n9414), .S(n6644), .Z(
        n4674) );
  MUX2_X2 U14182 ( .A(pipeline_regfile_data[508]), .B(n9415), .S(n6644), .Z(
        n4705) );
  MUX2_X2 U14183 ( .A(pipeline_regfile_data[505]), .B(n9418), .S(n6644), .Z(
        n4798) );
  MUX2_X2 U14184 ( .A(pipeline_regfile_data[503]), .B(n13005), .S(n6644), .Z(
        n4860) );
  MUX2_X2 U14185 ( .A(pipeline_regfile_data[502]), .B(n13006), .S(n6644), .Z(
        n4891) );
  MUX2_X2 U14186 ( .A(pipeline_regfile_data[501]), .B(n13007), .S(n6644), .Z(
        n4922) );
  MUX2_X2 U14187 ( .A(pipeline_regfile_data[499]), .B(n13009), .S(n6644), .Z(
        n4984) );
  MUX2_X2 U14188 ( .A(pipeline_regfile_data[498]), .B(n13010), .S(n6644), .Z(
        n5015) );
  MUX2_X2 U14189 ( .A(pipeline_regfile_data[496]), .B(n13012), .S(n6644), .Z(
        n5077) );
  MUX2_X2 U14190 ( .A(pipeline_regfile_data[495]), .B(n9420), .S(n6644), .Z(
        n5108) );
  MUX2_X2 U14191 ( .A(pipeline_regfile_data[494]), .B(n9421), .S(n6644), .Z(
        n5139) );
  MUX2_X2 U14192 ( .A(pipeline_regfile_data[490]), .B(n9427), .S(n6644), .Z(
        n5263) );
  MUX2_X2 U14193 ( .A(pipeline_regfile_data[489]), .B(n9429), .S(n6644), .Z(
        n5294) );
  MUX2_X2 U14194 ( .A(pipeline_regfile_data[488]), .B(n9431), .S(n6644), .Z(
        n5325) );
  MUX2_X2 U14195 ( .A(pipeline_regfile_data[487]), .B(n13021), .S(n6644), .Z(
        n5356) );
  MUX2_X2 U14196 ( .A(pipeline_regfile_data[485]), .B(n9433), .S(n6644), .Z(
        n5418) );
  MUX2_X2 U14197 ( .A(pipeline_regfile_data[484]), .B(n9434), .S(n6644), .Z(
        n5449) );
  MUX2_X2 U14198 ( .A(pipeline_regfile_data[480]), .B(n9438), .S(n6644), .Z(
        n5573) );
  MUX2_X2 U14199 ( .A(pipeline_regfile_data[479]), .B(n12997), .S(n6645), .Z(
        n4611) );
  MUX2_X2 U14200 ( .A(pipeline_regfile_data[478]), .B(n12998), .S(n6645), .Z(
        n4642) );
  MUX2_X2 U14201 ( .A(pipeline_regfile_data[477]), .B(n12999), .S(n6645), .Z(
        n4673) );
  MUX2_X2 U14202 ( .A(pipeline_regfile_data[476]), .B(n13000), .S(n6645), .Z(
        n4704) );
  MUX2_X2 U14203 ( .A(pipeline_regfile_data[473]), .B(n13003), .S(n6645), .Z(
        n4797) );
  MUX2_X2 U14204 ( .A(pipeline_regfile_data[471]), .B(n13005), .S(n6645), .Z(
        n4859) );
  MUX2_X2 U14205 ( .A(pipeline_regfile_data[470]), .B(n13006), .S(n6645), .Z(
        n4890) );
  MUX2_X2 U14206 ( .A(pipeline_regfile_data[469]), .B(n13007), .S(n6645), .Z(
        n4921) );
  MUX2_X2 U14207 ( .A(pipeline_regfile_data[467]), .B(n13009), .S(n6645), .Z(
        n4983) );
  MUX2_X2 U14208 ( .A(pipeline_regfile_data[466]), .B(n13010), .S(n6645), .Z(
        n5014) );
  MUX2_X2 U14209 ( .A(pipeline_regfile_data[464]), .B(n13012), .S(n6645), .Z(
        n5076) );
  MUX2_X2 U14210 ( .A(pipeline_regfile_data[463]), .B(n13013), .S(n6645), .Z(
        n5107) );
  MUX2_X2 U14211 ( .A(pipeline_regfile_data[462]), .B(n13014), .S(n6645), .Z(
        n5138) );
  MUX2_X2 U14212 ( .A(pipeline_regfile_data[458]), .B(n13018), .S(n6645), .Z(
        n5262) );
  MUX2_X2 U14213 ( .A(pipeline_regfile_data[457]), .B(n13019), .S(n6645), .Z(
        n5293) );
  MUX2_X2 U14214 ( .A(pipeline_regfile_data[456]), .B(n13020), .S(n6645), .Z(
        n5324) );
  MUX2_X2 U14215 ( .A(pipeline_regfile_data[455]), .B(n13021), .S(n6645), .Z(
        n5355) );
  MUX2_X2 U14216 ( .A(pipeline_regfile_data[453]), .B(n13023), .S(n6645), .Z(
        n5417) );
  MUX2_X2 U14217 ( .A(pipeline_regfile_data[452]), .B(n13024), .S(n6645), .Z(
        n5448) );
  MUX2_X2 U14218 ( .A(pipeline_regfile_data[451]), .B(n13025), .S(n6645), .Z(
        n5479) );
  MUX2_X2 U14219 ( .A(pipeline_regfile_data[448]), .B(n13028), .S(n6645), .Z(
        n5572) );
  MUX2_X2 U14220 ( .A(pipeline_regfile_data[447]), .B(n9412), .S(n6646), .Z(
        n4610) );
  MUX2_X2 U14221 ( .A(pipeline_regfile_data[446]), .B(n9413), .S(n6646), .Z(
        n4641) );
  MUX2_X2 U14222 ( .A(pipeline_regfile_data[445]), .B(n9414), .S(n6646), .Z(
        n4672) );
  MUX2_X2 U14223 ( .A(pipeline_regfile_data[444]), .B(n9415), .S(n6646), .Z(
        n4703) );
  MUX2_X2 U14224 ( .A(pipeline_regfile_data[441]), .B(n9418), .S(n6646), .Z(
        n4796) );
  MUX2_X2 U14225 ( .A(pipeline_regfile_data[439]), .B(n13005), .S(n6646), .Z(
        n4858) );
  MUX2_X2 U14226 ( .A(pipeline_regfile_data[438]), .B(n13006), .S(n6646), .Z(
        n4889) );
  MUX2_X2 U14227 ( .A(pipeline_regfile_data[437]), .B(n13007), .S(n6646), .Z(
        n4920) );
  MUX2_X2 U14228 ( .A(pipeline_regfile_data[435]), .B(n13009), .S(n6646), .Z(
        n4982) );
  MUX2_X2 U14229 ( .A(pipeline_regfile_data[434]), .B(n13010), .S(n6646), .Z(
        n5013) );
  MUX2_X2 U14230 ( .A(pipeline_regfile_data[432]), .B(n13012), .S(n6646), .Z(
        n5075) );
  MUX2_X2 U14231 ( .A(pipeline_regfile_data[431]), .B(n9420), .S(n6646), .Z(
        n5106) );
  MUX2_X2 U14232 ( .A(pipeline_regfile_data[430]), .B(n9421), .S(n6646), .Z(
        n5137) );
  MUX2_X2 U14233 ( .A(pipeline_regfile_data[426]), .B(n9426), .S(n6646), .Z(
        n5261) );
  MUX2_X2 U14234 ( .A(pipeline_regfile_data[425]), .B(n9428), .S(n6646), .Z(
        n5292) );
  MUX2_X2 U14235 ( .A(pipeline_regfile_data[424]), .B(n9430), .S(n6646), .Z(
        n5323) );
  MUX2_X2 U14236 ( .A(pipeline_regfile_data[423]), .B(n13021), .S(n6646), .Z(
        n5354) );
  MUX2_X2 U14237 ( .A(pipeline_regfile_data[421]), .B(n9433), .S(n6646), .Z(
        n5416) );
  MUX2_X2 U14238 ( .A(pipeline_regfile_data[420]), .B(n9434), .S(n6646), .Z(
        n5447) );
  MUX2_X2 U14239 ( .A(pipeline_regfile_data[419]), .B(n9435), .S(n6646), .Z(
        n5478) );
  MUX2_X2 U14240 ( .A(pipeline_regfile_data[416]), .B(n9438), .S(n6646), .Z(
        n5571) );
  MUX2_X2 U14241 ( .A(pipeline_regfile_data[415]), .B(n12997), .S(n6647), .Z(
        n4609) );
  MUX2_X2 U14242 ( .A(pipeline_regfile_data[414]), .B(n12998), .S(n6647), .Z(
        n4640) );
  MUX2_X2 U14243 ( .A(pipeline_regfile_data[413]), .B(n12999), .S(n6647), .Z(
        n4671) );
  MUX2_X2 U14244 ( .A(pipeline_regfile_data[412]), .B(n13000), .S(n6647), .Z(
        n4702) );
  MUX2_X2 U14245 ( .A(pipeline_regfile_data[409]), .B(n13003), .S(n6647), .Z(
        n4795) );
  MUX2_X2 U14246 ( .A(pipeline_regfile_data[407]), .B(n13005), .S(n6647), .Z(
        n4857) );
  MUX2_X2 U14247 ( .A(pipeline_regfile_data[406]), .B(n13006), .S(n6647), .Z(
        n4888) );
  MUX2_X2 U14248 ( .A(pipeline_regfile_data[405]), .B(n13007), .S(n6647), .Z(
        n4919) );
  MUX2_X2 U14249 ( .A(pipeline_regfile_data[403]), .B(n13009), .S(n6647), .Z(
        n4981) );
  MUX2_X2 U14250 ( .A(pipeline_regfile_data[402]), .B(n13010), .S(n6647), .Z(
        n5012) );
  MUX2_X2 U14251 ( .A(pipeline_regfile_data[400]), .B(n13012), .S(n6647), .Z(
        n5074) );
  MUX2_X2 U14252 ( .A(pipeline_regfile_data[399]), .B(n13013), .S(n6647), .Z(
        n5105) );
  MUX2_X2 U14253 ( .A(pipeline_regfile_data[398]), .B(n13014), .S(n6647), .Z(
        n5136) );
  MUX2_X2 U14254 ( .A(pipeline_regfile_data[394]), .B(n9427), .S(n6647), .Z(
        n5260) );
  MUX2_X2 U14255 ( .A(pipeline_regfile_data[393]), .B(n9429), .S(n6647), .Z(
        n5291) );
  MUX2_X2 U14256 ( .A(pipeline_regfile_data[392]), .B(n9431), .S(n6647), .Z(
        n5322) );
  MUX2_X2 U14257 ( .A(pipeline_regfile_data[391]), .B(n13021), .S(n6647), .Z(
        n5353) );
  MUX2_X2 U14258 ( .A(pipeline_regfile_data[389]), .B(n13023), .S(n6647), .Z(
        n5415) );
  MUX2_X2 U14259 ( .A(pipeline_regfile_data[388]), .B(n13024), .S(n6647), .Z(
        n5446) );
  MUX2_X2 U14260 ( .A(pipeline_regfile_data[387]), .B(n13025), .S(n6647), .Z(
        n5477) );
  MUX2_X2 U14261 ( .A(pipeline_regfile_data[384]), .B(n13028), .S(n6647), .Z(
        n5570) );
  MUX2_X2 U14262 ( .A(pipeline_regfile_data[383]), .B(n9412), .S(n6648), .Z(
        n4608) );
  MUX2_X2 U14263 ( .A(pipeline_regfile_data[382]), .B(n9413), .S(n6648), .Z(
        n4639) );
  MUX2_X2 U14264 ( .A(pipeline_regfile_data[381]), .B(n9414), .S(n6648), .Z(
        n4670) );
  MUX2_X2 U14265 ( .A(pipeline_regfile_data[380]), .B(n9415), .S(n6648), .Z(
        n4701) );
  MUX2_X2 U14266 ( .A(pipeline_regfile_data[377]), .B(n9418), .S(n6648), .Z(
        n4794) );
  MUX2_X2 U14267 ( .A(pipeline_regfile_data[376]), .B(n9419), .S(n6648), .Z(
        n4825) );
  MUX2_X2 U14268 ( .A(pipeline_regfile_data[375]), .B(n13005), .S(n6648), .Z(
        n4856) );
  MUX2_X2 U14269 ( .A(pipeline_regfile_data[374]), .B(n13006), .S(n6648), .Z(
        n4887) );
  MUX2_X2 U14270 ( .A(pipeline_regfile_data[373]), .B(n13007), .S(n6648), .Z(
        n4918) );
  MUX2_X2 U14271 ( .A(pipeline_regfile_data[372]), .B(n13008), .S(n6648), .Z(
        n4949) );
  MUX2_X2 U14272 ( .A(pipeline_regfile_data[371]), .B(n13009), .S(n6648), .Z(
        n4980) );
  MUX2_X2 U14273 ( .A(pipeline_regfile_data[370]), .B(n13010), .S(n6648), .Z(
        n5011) );
  MUX2_X2 U14274 ( .A(pipeline_regfile_data[368]), .B(n13012), .S(n6648), .Z(
        n5073) );
  MUX2_X2 U14275 ( .A(pipeline_regfile_data[367]), .B(n9420), .S(n6648), .Z(
        n5104) );
  MUX2_X2 U14276 ( .A(pipeline_regfile_data[366]), .B(n9421), .S(n6648), .Z(
        n5135) );
  MUX2_X2 U14277 ( .A(pipeline_regfile_data[365]), .B(n9422), .S(n6648), .Z(
        n5166) );
  MUX2_X2 U14278 ( .A(pipeline_regfile_data[363]), .B(n13017), .S(n6648), .Z(
        n5228) );
  MUX2_X2 U14279 ( .A(pipeline_regfile_data[362]), .B(n13018), .S(n6648), .Z(
        n5259) );
  MUX2_X2 U14280 ( .A(pipeline_regfile_data[361]), .B(n13019), .S(n6648), .Z(
        n5290) );
  MUX2_X2 U14281 ( .A(pipeline_regfile_data[360]), .B(n13020), .S(n6648), .Z(
        n5321) );
  MUX2_X2 U14282 ( .A(pipeline_regfile_data[359]), .B(n13021), .S(n6648), .Z(
        n5352) );
  MUX2_X2 U14283 ( .A(pipeline_regfile_data[357]), .B(n9433), .S(n6648), .Z(
        n5414) );
  MUX2_X2 U14284 ( .A(pipeline_regfile_data[355]), .B(n9435), .S(n6648), .Z(
        n5476) );
  MUX2_X2 U14285 ( .A(pipeline_regfile_data[352]), .B(n9438), .S(n6648), .Z(
        n5569) );
  MUX2_X2 U14286 ( .A(pipeline_regfile_data[351]), .B(n12997), .S(n6653), .Z(
        n4607) );
  MUX2_X2 U14287 ( .A(pipeline_regfile_data[350]), .B(n12998), .S(n6653), .Z(
        n4638) );
  MUX2_X2 U14288 ( .A(pipeline_regfile_data[349]), .B(n12999), .S(n6653), .Z(
        n4669) );
  MUX2_X2 U14289 ( .A(pipeline_regfile_data[348]), .B(n13000), .S(n6653), .Z(
        n4700) );
  MUX2_X2 U14290 ( .A(pipeline_regfile_data[347]), .B(n13001), .S(n6653), .Z(
        n4731) );
  MUX2_X2 U14291 ( .A(pipeline_regfile_data[345]), .B(n13003), .S(n6653), .Z(
        n4793) );
  MUX2_X2 U14292 ( .A(pipeline_regfile_data[344]), .B(n13004), .S(n6653), .Z(
        n4824) );
  MUX2_X2 U14293 ( .A(pipeline_regfile_data[343]), .B(n13005), .S(n6653), .Z(
        n4855) );
  MUX2_X2 U14294 ( .A(pipeline_regfile_data[342]), .B(n13006), .S(n6653), .Z(
        n4886) );
  MUX2_X2 U14295 ( .A(pipeline_regfile_data[341]), .B(n13007), .S(n6653), .Z(
        n4917) );
  MUX2_X2 U14296 ( .A(pipeline_regfile_data[340]), .B(n13008), .S(n6653), .Z(
        n4948) );
  MUX2_X2 U14297 ( .A(pipeline_regfile_data[339]), .B(n13009), .S(n6653), .Z(
        n4979) );
  MUX2_X2 U14298 ( .A(pipeline_regfile_data[338]), .B(n13010), .S(n6653), .Z(
        n5010) );
  MUX2_X2 U14299 ( .A(pipeline_regfile_data[337]), .B(n13011), .S(n6653), .Z(
        n5041) );
  MUX2_X2 U14300 ( .A(pipeline_regfile_data[336]), .B(n13012), .S(n6653), .Z(
        n5072) );
  MUX2_X2 U14301 ( .A(pipeline_regfile_data[335]), .B(n13013), .S(n6653), .Z(
        n5103) );
  MUX2_X2 U14302 ( .A(pipeline_regfile_data[334]), .B(n13014), .S(n6653), .Z(
        n5134) );
  MUX2_X2 U14303 ( .A(pipeline_regfile_data[333]), .B(n13015), .S(n6653), .Z(
        n5165) );
  MUX2_X2 U14304 ( .A(pipeline_regfile_data[331]), .B(n9424), .S(n6653), .Z(
        n5227) );
  MUX2_X2 U14305 ( .A(pipeline_regfile_data[330]), .B(n9426), .S(n6653), .Z(
        n5258) );
  MUX2_X2 U14306 ( .A(pipeline_regfile_data[329]), .B(n9428), .S(n6653), .Z(
        n5289) );
  MUX2_X2 U14307 ( .A(pipeline_regfile_data[328]), .B(n9430), .S(n6653), .Z(
        n5320) );
  MUX2_X2 U14308 ( .A(pipeline_regfile_data[327]), .B(n13021), .S(n6653), .Z(
        n5351) );
  MUX2_X2 U14309 ( .A(pipeline_regfile_data[325]), .B(n13023), .S(n6653), .Z(
        n5413) );
  MUX2_X2 U14310 ( .A(pipeline_regfile_data[323]), .B(n13025), .S(n6653), .Z(
        n5475) );
  MUX2_X2 U14311 ( .A(pipeline_regfile_data[320]), .B(n13028), .S(n6653), .Z(
        n5568) );
  MUX2_X2 U14312 ( .A(pipeline_regfile_data[319]), .B(n9412), .S(n6656), .Z(
        n4606) );
  MUX2_X2 U14313 ( .A(pipeline_regfile_data[318]), .B(n9413), .S(n6656), .Z(
        n4637) );
  MUX2_X2 U14314 ( .A(pipeline_regfile_data[317]), .B(n9414), .S(n6656), .Z(
        n4668) );
  MUX2_X2 U14315 ( .A(pipeline_regfile_data[316]), .B(n9415), .S(n6656), .Z(
        n4699) );
  MUX2_X2 U14316 ( .A(pipeline_regfile_data[315]), .B(n9416), .S(n6656), .Z(
        n4730) );
  MUX2_X2 U14317 ( .A(pipeline_regfile_data[314]), .B(n9417), .S(n6656), .Z(
        n4761) );
  MUX2_X2 U14318 ( .A(pipeline_regfile_data[313]), .B(n9418), .S(n6656), .Z(
        n4792) );
  MUX2_X2 U14319 ( .A(pipeline_regfile_data[312]), .B(n9419), .S(n6656), .Z(
        n4823) );
  MUX2_X2 U14320 ( .A(pipeline_regfile_data[311]), .B(n13005), .S(n6656), .Z(
        n4854) );
  MUX2_X2 U14321 ( .A(pipeline_regfile_data[310]), .B(n13006), .S(n6656), .Z(
        n4885) );
  MUX2_X2 U14322 ( .A(pipeline_regfile_data[309]), .B(n13007), .S(n6656), .Z(
        n4916) );
  MUX2_X2 U14323 ( .A(pipeline_regfile_data[308]), .B(n13008), .S(n6656), .Z(
        n4947) );
  MUX2_X2 U14324 ( .A(pipeline_regfile_data[307]), .B(n13009), .S(n6656), .Z(
        n4978) );
  MUX2_X2 U14325 ( .A(pipeline_regfile_data[306]), .B(n13010), .S(n6656), .Z(
        n5009) );
  MUX2_X2 U14326 ( .A(pipeline_regfile_data[305]), .B(n13011), .S(n6656), .Z(
        n5040) );
  MUX2_X2 U14327 ( .A(pipeline_regfile_data[304]), .B(n13012), .S(n6656), .Z(
        n5071) );
  MUX2_X2 U14328 ( .A(pipeline_regfile_data[303]), .B(n9420), .S(n6656), .Z(
        n5102) );
  MUX2_X2 U14329 ( .A(pipeline_regfile_data[302]), .B(n9421), .S(n6656), .Z(
        n5133) );
  MUX2_X2 U14330 ( .A(pipeline_regfile_data[301]), .B(n9422), .S(n6656), .Z(
        n5164) );
  MUX2_X2 U14331 ( .A(pipeline_regfile_data[299]), .B(n9425), .S(n6656), .Z(
        n5226) );
  MUX2_X2 U14332 ( .A(pipeline_regfile_data[298]), .B(n9427), .S(n6656), .Z(
        n5257) );
  MUX2_X2 U14333 ( .A(pipeline_regfile_data[297]), .B(n9429), .S(n6656), .Z(
        n5288) );
  MUX2_X2 U14334 ( .A(pipeline_regfile_data[296]), .B(n9431), .S(n6656), .Z(
        n5319) );
  MUX2_X2 U14335 ( .A(pipeline_regfile_data[295]), .B(n13021), .S(n6656), .Z(
        n5350) );
  MUX2_X2 U14336 ( .A(pipeline_regfile_data[294]), .B(n9432), .S(n6656), .Z(
        n5381) );
  MUX2_X2 U14337 ( .A(pipeline_regfile_data[293]), .B(n9433), .S(n6656), .Z(
        n5412) );
  MUX2_X2 U14338 ( .A(pipeline_regfile_data[292]), .B(n9434), .S(n6656), .Z(
        n5443) );
  MUX2_X2 U14339 ( .A(pipeline_regfile_data[291]), .B(n9435), .S(n6656), .Z(
        n5474) );
  MUX2_X2 U14340 ( .A(pipeline_regfile_data[288]), .B(n9438), .S(n6656), .Z(
        n5567) );
  MUX2_X2 U14341 ( .A(pipeline_regfile_data[287]), .B(n12997), .S(n6657), .Z(
        n4605) );
  MUX2_X2 U14342 ( .A(pipeline_regfile_data[286]), .B(n12998), .S(n6657), .Z(
        n4636) );
  MUX2_X2 U14343 ( .A(pipeline_regfile_data[285]), .B(n12999), .S(n6657), .Z(
        n4667) );
  MUX2_X2 U14344 ( .A(pipeline_regfile_data[284]), .B(n13000), .S(n6657), .Z(
        n4698) );
  MUX2_X2 U14345 ( .A(pipeline_regfile_data[283]), .B(n13001), .S(n6657), .Z(
        n4729) );
  MUX2_X2 U14346 ( .A(pipeline_regfile_data[282]), .B(n13002), .S(n6657), .Z(
        n4760) );
  MUX2_X2 U14347 ( .A(pipeline_regfile_data[281]), .B(n13003), .S(n6657), .Z(
        n4791) );
  MUX2_X2 U14348 ( .A(pipeline_regfile_data[280]), .B(n13004), .S(n6657), .Z(
        n4822) );
  MUX2_X2 U14349 ( .A(pipeline_regfile_data[279]), .B(n13005), .S(n6657), .Z(
        n4853) );
  MUX2_X2 U14350 ( .A(pipeline_regfile_data[278]), .B(n13006), .S(n6657), .Z(
        n4884) );
  MUX2_X2 U14351 ( .A(pipeline_regfile_data[277]), .B(n13007), .S(n6657), .Z(
        n4915) );
  MUX2_X2 U14352 ( .A(pipeline_regfile_data[276]), .B(n13008), .S(n6657), .Z(
        n4946) );
  MUX2_X2 U14353 ( .A(pipeline_regfile_data[275]), .B(n13009), .S(n6657), .Z(
        n4977) );
  MUX2_X2 U14354 ( .A(pipeline_regfile_data[274]), .B(n13010), .S(n6657), .Z(
        n5008) );
  MUX2_X2 U14355 ( .A(pipeline_regfile_data[273]), .B(n13011), .S(n6657), .Z(
        n5039) );
  MUX2_X2 U14356 ( .A(pipeline_regfile_data[272]), .B(n13012), .S(n6657), .Z(
        n5070) );
  MUX2_X2 U14357 ( .A(pipeline_regfile_data[271]), .B(n13013), .S(n6657), .Z(
        n5101) );
  MUX2_X2 U14358 ( .A(pipeline_regfile_data[270]), .B(n13014), .S(n6657), .Z(
        n5132) );
  MUX2_X2 U14359 ( .A(pipeline_regfile_data[269]), .B(n13015), .S(n6657), .Z(
        n5163) );
  MUX2_X2 U14360 ( .A(pipeline_regfile_data[267]), .B(n13017), .S(n6657), .Z(
        n5225) );
  MUX2_X2 U14361 ( .A(pipeline_regfile_data[266]), .B(n13018), .S(n6657), .Z(
        n5256) );
  MUX2_X2 U14362 ( .A(pipeline_regfile_data[265]), .B(n13019), .S(n6657), .Z(
        n5287) );
  MUX2_X2 U14363 ( .A(pipeline_regfile_data[264]), .B(n13020), .S(n6657), .Z(
        n5318) );
  MUX2_X2 U14364 ( .A(pipeline_regfile_data[263]), .B(n13021), .S(n6657), .Z(
        n5349) );
  MUX2_X2 U14365 ( .A(pipeline_regfile_data[262]), .B(n13022), .S(n6657), .Z(
        n5380) );
  MUX2_X2 U14366 ( .A(pipeline_regfile_data[261]), .B(n13023), .S(n6657), .Z(
        n5411) );
  MUX2_X2 U14367 ( .A(pipeline_regfile_data[260]), .B(n13024), .S(n6657), .Z(
        n5442) );
  MUX2_X2 U14368 ( .A(pipeline_regfile_data[259]), .B(n13025), .S(n6657), .Z(
        n5473) );
  MUX2_X2 U14369 ( .A(pipeline_regfile_data[258]), .B(n13026), .S(n6657), .Z(
        n5504) );
  MUX2_X2 U14370 ( .A(pipeline_regfile_data[256]), .B(n13028), .S(n6657), .Z(
        n5566) );
  MUX2_X2 U14371 ( .A(pipeline_regfile_data[255]), .B(n9412), .S(n6649), .Z(
        n4604) );
  MUX2_X2 U14372 ( .A(pipeline_regfile_data[254]), .B(n9413), .S(n6649), .Z(
        n4635) );
  MUX2_X2 U14373 ( .A(pipeline_regfile_data[253]), .B(n9414), .S(n6649), .Z(
        n4666) );
  MUX2_X2 U14374 ( .A(pipeline_regfile_data[252]), .B(n9415), .S(n6649), .Z(
        n4697) );
  MUX2_X2 U14375 ( .A(pipeline_regfile_data[251]), .B(n9416), .S(n6649), .Z(
        n4728) );
  MUX2_X2 U14376 ( .A(pipeline_regfile_data[249]), .B(n9418), .S(n6649), .Z(
        n4790) );
  MUX2_X2 U14377 ( .A(pipeline_regfile_data[247]), .B(n13005), .S(n6649), .Z(
        n4852) );
  MUX2_X2 U14378 ( .A(pipeline_regfile_data[246]), .B(n13006), .S(n6649), .Z(
        n4883) );
  MUX2_X2 U14379 ( .A(pipeline_regfile_data[245]), .B(n13007), .S(n6649), .Z(
        n4914) );
  MUX2_X2 U14380 ( .A(pipeline_regfile_data[243]), .B(n13009), .S(n6649), .Z(
        n4976) );
  MUX2_X2 U14381 ( .A(pipeline_regfile_data[242]), .B(n13010), .S(n6649), .Z(
        n5007) );
  MUX2_X2 U14382 ( .A(pipeline_regfile_data[240]), .B(n13012), .S(n6649), .Z(
        n5069) );
  MUX2_X2 U14383 ( .A(pipeline_regfile_data[239]), .B(n9420), .S(n6649), .Z(
        n5100) );
  MUX2_X2 U14384 ( .A(pipeline_regfile_data[238]), .B(n9421), .S(n6649), .Z(
        n5131) );
  MUX2_X2 U14385 ( .A(pipeline_regfile_data[237]), .B(n9422), .S(n6649), .Z(
        n5162) );
  MUX2_X2 U14386 ( .A(pipeline_regfile_data[235]), .B(n9424), .S(n6649), .Z(
        n5224) );
  MUX2_X2 U14387 ( .A(pipeline_regfile_data[234]), .B(n9426), .S(n6649), .Z(
        n5255) );
  MUX2_X2 U14388 ( .A(pipeline_regfile_data[233]), .B(n9428), .S(n6649), .Z(
        n5286) );
  MUX2_X2 U14389 ( .A(pipeline_regfile_data[232]), .B(n9430), .S(n6649), .Z(
        n5317) );
  MUX2_X2 U14390 ( .A(pipeline_regfile_data[231]), .B(n13021), .S(n6649), .Z(
        n5348) );
  MUX2_X2 U14391 ( .A(pipeline_regfile_data[229]), .B(n9433), .S(n6649), .Z(
        n5410) );
  MUX2_X2 U14392 ( .A(pipeline_regfile_data[228]), .B(n9434), .S(n6649), .Z(
        n5441) );
  MUX2_X2 U14393 ( .A(pipeline_regfile_data[227]), .B(n9435), .S(n6649), .Z(
        n5472) );
  MUX2_X2 U14394 ( .A(pipeline_regfile_data[224]), .B(n9438), .S(n6649), .Z(
        n5565) );
  MUX2_X2 U14395 ( .A(pipeline_regfile_data[223]), .B(n12997), .S(n6650), .Z(
        n4603) );
  MUX2_X2 U14396 ( .A(pipeline_regfile_data[222]), .B(n12998), .S(n6650), .Z(
        n4634) );
  MUX2_X2 U14397 ( .A(pipeline_regfile_data[221]), .B(n12999), .S(n6650), .Z(
        n4665) );
  MUX2_X2 U14398 ( .A(pipeline_regfile_data[220]), .B(n13000), .S(n6650), .Z(
        n4696) );
  MUX2_X2 U14399 ( .A(pipeline_regfile_data[219]), .B(n13001), .S(n6650), .Z(
        n4727) );
  MUX2_X2 U14400 ( .A(pipeline_regfile_data[217]), .B(n13003), .S(n6650), .Z(
        n4789) );
  MUX2_X2 U14401 ( .A(pipeline_regfile_data[215]), .B(n13005), .S(n6650), .Z(
        n4851) );
  MUX2_X2 U14402 ( .A(pipeline_regfile_data[214]), .B(n13006), .S(n6650), .Z(
        n4882) );
  MUX2_X2 U14403 ( .A(pipeline_regfile_data[213]), .B(n13007), .S(n6650), .Z(
        n4913) );
  MUX2_X2 U14404 ( .A(pipeline_regfile_data[211]), .B(n13009), .S(n6650), .Z(
        n4975) );
  MUX2_X2 U14405 ( .A(pipeline_regfile_data[210]), .B(n13010), .S(n6650), .Z(
        n5006) );
  MUX2_X2 U14406 ( .A(pipeline_regfile_data[208]), .B(n13012), .S(n6650), .Z(
        n5068) );
  MUX2_X2 U14407 ( .A(pipeline_regfile_data[207]), .B(n13013), .S(n6650), .Z(
        n5099) );
  MUX2_X2 U14408 ( .A(pipeline_regfile_data[206]), .B(n13014), .S(n6650), .Z(
        n5130) );
  MUX2_X2 U14409 ( .A(pipeline_regfile_data[205]), .B(n13015), .S(n6650), .Z(
        n5161) );
  MUX2_X2 U14410 ( .A(pipeline_regfile_data[203]), .B(n9425), .S(n6650), .Z(
        n5223) );
  MUX2_X2 U14411 ( .A(pipeline_regfile_data[202]), .B(n9427), .S(n6650), .Z(
        n5254) );
  MUX2_X2 U14412 ( .A(pipeline_regfile_data[201]), .B(n9429), .S(n6650), .Z(
        n5285) );
  MUX2_X2 U14413 ( .A(pipeline_regfile_data[200]), .B(n9431), .S(n6650), .Z(
        n5316) );
  MUX2_X2 U14414 ( .A(pipeline_regfile_data[199]), .B(n13021), .S(n6650), .Z(
        n5347) );
  MUX2_X2 U14415 ( .A(pipeline_regfile_data[197]), .B(n13023), .S(n6650), .Z(
        n5409) );
  MUX2_X2 U14416 ( .A(pipeline_regfile_data[196]), .B(n13024), .S(n6650), .Z(
        n5440) );
  MUX2_X2 U14417 ( .A(pipeline_regfile_data[195]), .B(n13025), .S(n6650), .Z(
        n5471) );
  MUX2_X2 U14418 ( .A(pipeline_regfile_data[192]), .B(n13028), .S(n6650), .Z(
        n5564) );
  MUX2_X2 U14419 ( .A(pipeline_regfile_data[191]), .B(n9412), .S(n6651), .Z(
        n4602) );
  MUX2_X2 U14420 ( .A(pipeline_regfile_data[190]), .B(n9413), .S(n6651), .Z(
        n4633) );
  MUX2_X2 U14421 ( .A(pipeline_regfile_data[189]), .B(n9414), .S(n6651), .Z(
        n4664) );
  MUX2_X2 U14422 ( .A(pipeline_regfile_data[188]), .B(n9415), .S(n6651), .Z(
        n4695) );
  MUX2_X2 U14423 ( .A(pipeline_regfile_data[187]), .B(n9416), .S(n6651), .Z(
        n4726) );
  MUX2_X2 U14424 ( .A(pipeline_regfile_data[185]), .B(n9418), .S(n6651), .Z(
        n4788) );
  MUX2_X2 U14425 ( .A(pipeline_regfile_data[183]), .B(n13005), .S(n6651), .Z(
        n4850) );
  MUX2_X2 U14426 ( .A(pipeline_regfile_data[182]), .B(n13006), .S(n6651), .Z(
        n4881) );
  MUX2_X2 U14427 ( .A(pipeline_regfile_data[181]), .B(n13007), .S(n6651), .Z(
        n4912) );
  MUX2_X2 U14428 ( .A(pipeline_regfile_data[179]), .B(n13009), .S(n6651), .Z(
        n4974) );
  MUX2_X2 U14429 ( .A(pipeline_regfile_data[178]), .B(n13010), .S(n6651), .Z(
        n5005) );
  MUX2_X2 U14430 ( .A(pipeline_regfile_data[176]), .B(n13012), .S(n6651), .Z(
        n5067) );
  MUX2_X2 U14431 ( .A(pipeline_regfile_data[175]), .B(n9420), .S(n6651), .Z(
        n5098) );
  MUX2_X2 U14432 ( .A(pipeline_regfile_data[174]), .B(n9421), .S(n6651), .Z(
        n5129) );
  MUX2_X2 U14433 ( .A(pipeline_regfile_data[173]), .B(n9422), .S(n6651), .Z(
        n5160) );
  MUX2_X2 U14434 ( .A(pipeline_regfile_data[171]), .B(n13017), .S(n6651), .Z(
        n5222) );
  MUX2_X2 U14435 ( .A(pipeline_regfile_data[170]), .B(n13018), .S(n6651), .Z(
        n5253) );
  MUX2_X2 U14436 ( .A(pipeline_regfile_data[169]), .B(n13019), .S(n6651), .Z(
        n5284) );
  MUX2_X2 U14437 ( .A(pipeline_regfile_data[168]), .B(n13020), .S(n6651), .Z(
        n5315) );
  MUX2_X2 U14438 ( .A(pipeline_regfile_data[167]), .B(n13021), .S(n6651), .Z(
        n5346) );
  MUX2_X2 U14439 ( .A(pipeline_regfile_data[165]), .B(n9433), .S(n6651), .Z(
        n5408) );
  MUX2_X2 U14440 ( .A(pipeline_regfile_data[164]), .B(n9434), .S(n6651), .Z(
        n5439) );
  MUX2_X2 U14441 ( .A(pipeline_regfile_data[163]), .B(n9435), .S(n6651), .Z(
        n5470) );
  MUX2_X2 U14442 ( .A(pipeline_regfile_data[160]), .B(n9438), .S(n6651), .Z(
        n5563) );
  MUX2_X2 U14443 ( .A(pipeline_regfile_data[159]), .B(n12997), .S(n6652), .Z(
        n4601) );
  MUX2_X2 U14444 ( .A(pipeline_regfile_data[158]), .B(n12998), .S(n6652), .Z(
        n4632) );
  MUX2_X2 U14445 ( .A(pipeline_regfile_data[157]), .B(n12999), .S(n6652), .Z(
        n4663) );
  MUX2_X2 U14446 ( .A(pipeline_regfile_data[156]), .B(n13000), .S(n6652), .Z(
        n4694) );
  MUX2_X2 U14447 ( .A(pipeline_regfile_data[155]), .B(n13001), .S(n6652), .Z(
        n4725) );
  MUX2_X2 U14448 ( .A(pipeline_regfile_data[153]), .B(n13003), .S(n6652), .Z(
        n4787) );
  MUX2_X2 U14449 ( .A(pipeline_regfile_data[151]), .B(n13005), .S(n6652), .Z(
        n4849) );
  MUX2_X2 U14450 ( .A(pipeline_regfile_data[150]), .B(n13006), .S(n6652), .Z(
        n4880) );
  MUX2_X2 U14451 ( .A(pipeline_regfile_data[149]), .B(n13007), .S(n6652), .Z(
        n4911) );
  MUX2_X2 U14452 ( .A(pipeline_regfile_data[147]), .B(n13009), .S(n6652), .Z(
        n4973) );
  MUX2_X2 U14453 ( .A(pipeline_regfile_data[146]), .B(n13010), .S(n6652), .Z(
        n5004) );
  MUX2_X2 U14454 ( .A(pipeline_regfile_data[144]), .B(n13012), .S(n6652), .Z(
        n5066) );
  MUX2_X2 U14455 ( .A(pipeline_regfile_data[143]), .B(n13013), .S(n6652), .Z(
        n5097) );
  MUX2_X2 U14456 ( .A(pipeline_regfile_data[142]), .B(n13014), .S(n6652), .Z(
        n5128) );
  MUX2_X2 U14457 ( .A(pipeline_regfile_data[141]), .B(n13015), .S(n6652), .Z(
        n5159) );
  MUX2_X2 U14458 ( .A(pipeline_regfile_data[139]), .B(n9424), .S(n6652), .Z(
        n5221) );
  MUX2_X2 U14459 ( .A(pipeline_regfile_data[138]), .B(n9426), .S(n6652), .Z(
        n5252) );
  MUX2_X2 U14460 ( .A(pipeline_regfile_data[137]), .B(n9428), .S(n6652), .Z(
        n5283) );
  MUX2_X2 U14461 ( .A(pipeline_regfile_data[136]), .B(n9430), .S(n6652), .Z(
        n5314) );
  MUX2_X2 U14462 ( .A(pipeline_regfile_data[135]), .B(n13021), .S(n6652), .Z(
        n5345) );
  MUX2_X2 U14463 ( .A(pipeline_regfile_data[133]), .B(n13023), .S(n6652), .Z(
        n5407) );
  MUX2_X2 U14464 ( .A(pipeline_regfile_data[132]), .B(n13024), .S(n6652), .Z(
        n5438) );
  MUX2_X2 U14465 ( .A(pipeline_regfile_data[131]), .B(n13025), .S(n6652), .Z(
        n5469) );
  MUX2_X2 U14466 ( .A(pipeline_regfile_data[128]), .B(n13028), .S(n6652), .Z(
        n5562) );
  MUX2_X2 U14467 ( .A(pipeline_regfile_data[127]), .B(n9412), .S(n6654), .Z(
        n4600) );
  MUX2_X2 U14468 ( .A(pipeline_regfile_data[126]), .B(n9413), .S(n6654), .Z(
        n4631) );
  MUX2_X2 U14469 ( .A(pipeline_regfile_data[125]), .B(n9414), .S(n6654), .Z(
        n4662) );
  MUX2_X2 U14470 ( .A(pipeline_regfile_data[124]), .B(n9415), .S(n6654), .Z(
        n4693) );
  MUX2_X2 U14471 ( .A(pipeline_regfile_data[123]), .B(n9416), .S(n6654), .Z(
        n4724) );
  MUX2_X2 U14472 ( .A(pipeline_regfile_data[121]), .B(n9418), .S(n6654), .Z(
        n4786) );
  MUX2_X2 U14473 ( .A(pipeline_regfile_data[120]), .B(n9419), .S(n6654), .Z(
        n4817) );
  MUX2_X2 U14474 ( .A(pipeline_regfile_data[119]), .B(n13005), .S(n6654), .Z(
        n4848) );
  MUX2_X2 U14475 ( .A(pipeline_regfile_data[118]), .B(n13006), .S(n6654), .Z(
        n4879) );
  MUX2_X2 U14476 ( .A(pipeline_regfile_data[117]), .B(n13007), .S(n6654), .Z(
        n4910) );
  MUX2_X2 U14477 ( .A(pipeline_regfile_data[116]), .B(n13008), .S(n6654), .Z(
        n4941) );
  MUX2_X2 U14478 ( .A(pipeline_regfile_data[115]), .B(n13009), .S(n6654), .Z(
        n4972) );
  MUX2_X2 U14479 ( .A(pipeline_regfile_data[114]), .B(n13010), .S(n6654), .Z(
        n5003) );
  MUX2_X2 U14480 ( .A(pipeline_regfile_data[113]), .B(n13011), .S(n6654), .Z(
        n5034) );
  MUX2_X2 U14481 ( .A(pipeline_regfile_data[112]), .B(n13012), .S(n6654), .Z(
        n5065) );
  MUX2_X2 U14482 ( .A(pipeline_regfile_data[111]), .B(n9420), .S(n6654), .Z(
        n5096) );
  MUX2_X2 U14483 ( .A(pipeline_regfile_data[110]), .B(n9421), .S(n6654), .Z(
        n5127) );
  MUX2_X2 U14484 ( .A(pipeline_regfile_data[109]), .B(n9422), .S(n6654), .Z(
        n5158) );
  MUX2_X2 U14485 ( .A(pipeline_regfile_data[107]), .B(n9425), .S(n6654), .Z(
        n5220) );
  MUX2_X2 U14486 ( .A(pipeline_regfile_data[106]), .B(n9427), .S(n6654), .Z(
        n5251) );
  MUX2_X2 U14487 ( .A(pipeline_regfile_data[105]), .B(n9429), .S(n6654), .Z(
        n5282) );
  MUX2_X2 U14488 ( .A(pipeline_regfile_data[104]), .B(n9431), .S(n6654), .Z(
        n5313) );
  MUX2_X2 U14489 ( .A(pipeline_regfile_data[103]), .B(n13021), .S(n6654), .Z(
        n5344) );
  MUX2_X2 U14490 ( .A(pipeline_regfile_data[101]), .B(n9433), .S(n6654), .Z(
        n5406) );
  MUX2_X2 U14491 ( .A(pipeline_regfile_data[99]), .B(n9435), .S(n6654), .Z(
        n5468) );
  MUX2_X2 U14492 ( .A(pipeline_regfile_data[96]), .B(n9438), .S(n6654), .Z(
        n5561) );
  MUX2_X2 U14493 ( .A(pipeline_regfile_data[95]), .B(n12997), .S(n6655), .Z(
        n4599) );
  MUX2_X2 U14494 ( .A(pipeline_regfile_data[94]), .B(n12998), .S(n6655), .Z(
        n4630) );
  MUX2_X2 U14495 ( .A(pipeline_regfile_data[93]), .B(n12999), .S(n6655), .Z(
        n4661) );
  MUX2_X2 U14496 ( .A(pipeline_regfile_data[92]), .B(n13000), .S(n6655), .Z(
        n4692) );
  MUX2_X2 U14497 ( .A(pipeline_regfile_data[91]), .B(n13001), .S(n6655), .Z(
        n4723) );
  MUX2_X2 U14498 ( .A(pipeline_regfile_data[89]), .B(n13003), .S(n6655), .Z(
        n4785) );
  MUX2_X2 U14499 ( .A(pipeline_regfile_data[88]), .B(n13004), .S(n6655), .Z(
        n4816) );
  MUX2_X2 U14500 ( .A(pipeline_regfile_data[87]), .B(n13005), .S(n6655), .Z(
        n4847) );
  MUX2_X2 U14501 ( .A(pipeline_regfile_data[86]), .B(n13006), .S(n6655), .Z(
        n4878) );
  MUX2_X2 U14502 ( .A(pipeline_regfile_data[85]), .B(n13007), .S(n6655), .Z(
        n4909) );
  MUX2_X2 U14503 ( .A(pipeline_regfile_data[84]), .B(n13008), .S(n6655), .Z(
        n4940) );
  MUX2_X2 U14504 ( .A(pipeline_regfile_data[83]), .B(n13009), .S(n6655), .Z(
        n4971) );
  MUX2_X2 U14505 ( .A(pipeline_regfile_data[82]), .B(n13010), .S(n6655), .Z(
        n5002) );
  MUX2_X2 U14506 ( .A(pipeline_regfile_data[81]), .B(n13011), .S(n6655), .Z(
        n5033) );
  MUX2_X2 U14507 ( .A(pipeline_regfile_data[80]), .B(n13012), .S(n6655), .Z(
        n5064) );
  MUX2_X2 U14508 ( .A(pipeline_regfile_data[79]), .B(n13013), .S(n6655), .Z(
        n5095) );
  MUX2_X2 U14509 ( .A(pipeline_regfile_data[78]), .B(n13014), .S(n6655), .Z(
        n5126) );
  MUX2_X2 U14510 ( .A(pipeline_regfile_data[77]), .B(n13015), .S(n6655), .Z(
        n5157) );
  MUX2_X2 U14511 ( .A(pipeline_regfile_data[75]), .B(n13017), .S(n6655), .Z(
        n5219) );
  MUX2_X2 U14512 ( .A(pipeline_regfile_data[74]), .B(n13018), .S(n6655), .Z(
        n5250) );
  MUX2_X2 U14513 ( .A(pipeline_regfile_data[73]), .B(n13019), .S(n6655), .Z(
        n5281) );
  MUX2_X2 U14514 ( .A(pipeline_regfile_data[72]), .B(n13020), .S(n6655), .Z(
        n5312) );
  MUX2_X2 U14515 ( .A(pipeline_regfile_data[71]), .B(n13021), .S(n6655), .Z(
        n5343) );
  MUX2_X2 U14516 ( .A(pipeline_regfile_data[69]), .B(n13023), .S(n6655), .Z(
        n5405) );
  MUX2_X2 U14517 ( .A(pipeline_regfile_data[67]), .B(n13025), .S(n6655), .Z(
        n5467) );
  MUX2_X2 U14518 ( .A(pipeline_regfile_data[64]), .B(n13028), .S(n6655), .Z(
        n5560) );
  MUX2_X2 U14519 ( .A(pipeline_regfile_data[63]), .B(n9412), .S(n6658), .Z(
        n4598) );
  MUX2_X2 U14520 ( .A(pipeline_regfile_data[62]), .B(n9413), .S(n6658), .Z(
        n4629) );
  MUX2_X2 U14521 ( .A(pipeline_regfile_data[61]), .B(n9414), .S(n6658), .Z(
        n4660) );
  MUX2_X2 U14522 ( .A(pipeline_regfile_data[60]), .B(n9415), .S(n6658), .Z(
        n4691) );
  MUX2_X2 U14523 ( .A(pipeline_regfile_data[59]), .B(n9416), .S(n6658), .Z(
        n4722) );
  MUX2_X2 U14524 ( .A(pipeline_regfile_data[58]), .B(n9417), .S(n6658), .Z(
        n4753) );
  MUX2_X2 U14525 ( .A(pipeline_regfile_data[57]), .B(n9418), .S(n6658), .Z(
        n4784) );
  MUX2_X2 U14526 ( .A(pipeline_regfile_data[56]), .B(n9419), .S(n6658), .Z(
        n4815) );
  MUX2_X2 U14527 ( .A(pipeline_regfile_data[55]), .B(n13005), .S(n6658), .Z(
        n4846) );
  MUX2_X2 U14528 ( .A(pipeline_regfile_data[54]), .B(n13006), .S(n6658), .Z(
        n4877) );
  MUX2_X2 U14529 ( .A(pipeline_regfile_data[53]), .B(n13007), .S(n6658), .Z(
        n4908) );
  MUX2_X2 U14530 ( .A(pipeline_regfile_data[52]), .B(n13008), .S(n6658), .Z(
        n4939) );
  MUX2_X2 U14531 ( .A(pipeline_regfile_data[51]), .B(n13009), .S(n6658), .Z(
        n4970) );
  MUX2_X2 U14532 ( .A(pipeline_regfile_data[50]), .B(n13010), .S(n6658), .Z(
        n5001) );
  MUX2_X2 U14533 ( .A(pipeline_regfile_data[49]), .B(n13011), .S(n6658), .Z(
        n5032) );
  MUX2_X2 U14534 ( .A(pipeline_regfile_data[48]), .B(n13012), .S(n6658), .Z(
        n5063) );
  MUX2_X2 U14535 ( .A(pipeline_regfile_data[47]), .B(n9420), .S(n6658), .Z(
        n5094) );
  MUX2_X2 U14536 ( .A(pipeline_regfile_data[46]), .B(n9421), .S(n6658), .Z(
        n5125) );
  MUX2_X2 U14537 ( .A(pipeline_regfile_data[45]), .B(n9422), .S(n6658), .Z(
        n5156) );
  MUX2_X2 U14538 ( .A(pipeline_regfile_data[43]), .B(n9424), .S(n6658), .Z(
        n5218) );
  MUX2_X2 U14539 ( .A(pipeline_regfile_data[42]), .B(n9426), .S(n6658), .Z(
        n5249) );
  MUX2_X2 U14540 ( .A(pipeline_regfile_data[41]), .B(n9428), .S(n6658), .Z(
        n5280) );
  MUX2_X2 U14541 ( .A(pipeline_regfile_data[40]), .B(n9430), .S(n6658), .Z(
        n5311) );
  MUX2_X2 U14542 ( .A(pipeline_regfile_data[39]), .B(n13021), .S(n6658), .Z(
        n5342) );
  MUX2_X2 U14543 ( .A(pipeline_regfile_data[38]), .B(n9432), .S(n6658), .Z(
        n5373) );
  MUX2_X2 U14544 ( .A(pipeline_regfile_data[37]), .B(n9433), .S(n6658), .Z(
        n5404) );
  MUX2_X2 U14545 ( .A(pipeline_regfile_data[36]), .B(n9434), .S(n6658), .Z(
        n5435) );
  MUX2_X2 U14546 ( .A(pipeline_regfile_data[35]), .B(n9435), .S(n6658), .Z(
        n5466) );
  MUX2_X2 U14547 ( .A(pipeline_regfile_data[34]), .B(n9436), .S(n6658), .Z(
        n5497) );
  MUX2_X2 U14548 ( .A(pipeline_regfile_data[32]), .B(n9438), .S(n6658), .Z(
        n5559) );
  MUX2_X2 U14550 ( .A(n13029), .B(n9521), .S(pipeline_md_N21), .Z(n13030) );
  NAND2_X2 U14551 ( .A1(n13031), .A2(n13030), .ZN(n6249) );
  AOI221_X2 U14552 ( .B1(pipeline_md_N181), .B2(n9519), .C1(n6643), .C2(
        pipeline_md_N23), .A(n13034), .ZN(n13032) );
  INV_X4 U14553 ( .A(n13032), .ZN(n6248) );
  AOI221_X2 U14554 ( .B1(pipeline_md_N182), .B2(n9519), .C1(pipeline_md_N24), 
        .C2(n6643), .A(n13034), .ZN(n13033) );
  INV_X4 U14555 ( .A(n13033), .ZN(n6247) );
  AOI221_X2 U14556 ( .B1(pipeline_md_N183), .B2(n9519), .C1(n6643), .C2(
        pipeline_md_N25), .A(n13034), .ZN(n13035) );
  INV_X4 U14557 ( .A(n13035), .ZN(n6246) );
  OAI22_X2 U14558 ( .A1(n6715), .A2(n13037), .B1(n6814), .B2(n13036), .ZN(
        n13038) );
  AOI221_X2 U14559 ( .B1(pipeline_md_a[9]), .B2(n142), .C1(pipeline_md_a[8]), 
        .C2(n143), .A(n13038), .ZN(n13043) );
  OAI22_X2 U14560 ( .A1(n6715), .A2(n13040), .B1(n6814), .B2(n13039), .ZN(
        n13041) );
  AOI221_X2 U14561 ( .B1(pipeline_md_a[13]), .B2(n142), .C1(pipeline_md_a[12]), 
        .C2(n143), .A(n13041), .ZN(n13042) );
  MUX2_X2 U14562 ( .A(n13043), .B(n13042), .S(pipeline_md_N23), .Z(n13044) );
  INV_X4 U14563 ( .A(n13044), .ZN(n150) );
  OAI22_X2 U14564 ( .A1(n6715), .A2(n13046), .B1(n6814), .B2(n13045), .ZN(
        n13047) );
  AOI221_X2 U14565 ( .B1(pipeline_md_a[1]), .B2(n142), .C1(pipeline_md_a[0]), 
        .C2(n143), .A(n13047), .ZN(n13052) );
  OAI22_X2 U14566 ( .A1(n6715), .A2(n13049), .B1(n6814), .B2(n13048), .ZN(
        n13050) );
  AOI221_X2 U14567 ( .B1(pipeline_md_a[5]), .B2(n142), .C1(pipeline_md_a[4]), 
        .C2(n143), .A(n13050), .ZN(n13051) );
  MUX2_X2 U14568 ( .A(n13052), .B(n13051), .S(pipeline_md_N23), .Z(n13053) );
  INV_X4 U14569 ( .A(n13053), .ZN(n149) );
  OAI22_X2 U14570 ( .A1(n6715), .A2(n13055), .B1(n6814), .B2(n13054), .ZN(
        n13056) );
  AOI221_X2 U14571 ( .B1(pipeline_md_a[25]), .B2(n142), .C1(pipeline_md_a[24]), 
        .C2(n143), .A(n13056), .ZN(n13061) );
  OAI22_X2 U14572 ( .A1(n6715), .A2(n13058), .B1(n6814), .B2(n13057), .ZN(
        n13059) );
  AOI221_X2 U14573 ( .B1(pipeline_md_a[29]), .B2(n142), .C1(pipeline_md_a[28]), 
        .C2(n143), .A(n13059), .ZN(n13060) );
  MUX2_X2 U14574 ( .A(n13061), .B(n13060), .S(pipeline_md_N23), .Z(n13062) );
  INV_X4 U14575 ( .A(n13062), .ZN(n136) );
  OAI22_X2 U14576 ( .A1(n6715), .A2(n13064), .B1(n6814), .B2(n13063), .ZN(
        n13065) );
  AOI221_X2 U14577 ( .B1(pipeline_md_a[17]), .B2(n142), .C1(pipeline_md_a[16]), 
        .C2(n143), .A(n13065), .ZN(n13070) );
  OAI22_X2 U14578 ( .A1(n6715), .A2(n13067), .B1(n6814), .B2(n13066), .ZN(
        n13068) );
  AOI221_X2 U14579 ( .B1(pipeline_md_a[21]), .B2(n142), .C1(pipeline_md_a[20]), 
        .C2(n143), .A(n13068), .ZN(n13069) );
  MUX2_X2 U14580 ( .A(n13070), .B(n13069), .S(pipeline_md_N23), .Z(n13071) );
  INV_X4 U14581 ( .A(n13071), .ZN(n135) );
  MUX2_X2 U14582 ( .A(n13072), .B(pipeline_rs2_data_bypassed[10]), .S(n9522), 
        .Z(n6322) );
  MUX2_X2 U14583 ( .A(dmem_hwdata[2]), .B(pipeline_rs2_data_bypassed[2]), .S(
        n9523), .Z(n6330) );
  MUX2_X2 U14584 ( .A(n13073), .B(pipeline_rs2_data_bypassed[11]), .S(n9524), 
        .Z(n6321) );
  MUX2_X2 U14585 ( .A(dmem_hwdata[3]), .B(n6987), .S(n9522), .Z(n6329) );
  MUX2_X2 U14586 ( .A(n13074), .B(pipeline_rs2_data_bypassed[12]), .S(n9523), 
        .Z(n6320) );
  MUX2_X2 U14587 ( .A(dmem_hwdata[4]), .B(n7004), .S(n9524), .Z(n6328) );
  MUX2_X2 U14588 ( .A(n13075), .B(pipeline_rs2_data_bypassed[13]), .S(n9524), 
        .Z(n6319) );
  MUX2_X2 U14589 ( .A(dmem_hwdata[5]), .B(pipeline_rs2_data_bypassed[5]), .S(
        n9522), .Z(n6327) );
  MUX2_X2 U14590 ( .A(n13076), .B(pipeline_rs2_data_bypassed[14]), .S(n9525), 
        .Z(n6318) );
  MUX2_X2 U14591 ( .A(dmem_hwdata[6]), .B(pipeline_rs2_data_bypassed[6]), .S(
        n9524), .Z(n6326) );
  MUX2_X2 U14592 ( .A(n13077), .B(pipeline_rs2_data_bypassed[15]), .S(n9522), 
        .Z(n6317) );
  MUX2_X2 U14593 ( .A(dmem_hwdata[7]), .B(pipeline_rs2_data_bypassed[7]), .S(
        n9525), .Z(n6325) );
  MUX2_X2 U14594 ( .A(dmem_hwdata[0]), .B(pipeline_rs2_data_bypassed[0]), .S(
        n9525), .Z(n6332) );
  MUX2_X2 U14595 ( .A(n13078), .B(pipeline_rs2_data_bypassed[16]), .S(n9522), 
        .Z(n6316) );
  MUX2_X2 U14596 ( .A(dmem_hwdata[1]), .B(pipeline_rs2_data_bypassed[1]), .S(
        n9523), .Z(n6331) );
  MUX2_X2 U14597 ( .A(n13079), .B(pipeline_rs2_data_bypassed[17]), .S(n9522), 
        .Z(n6315) );
  MUX2_X2 U14598 ( .A(n13080), .B(pipeline_rs2_data_bypassed[18]), .S(n9524), 
        .Z(n6314) );
  MUX2_X2 U14599 ( .A(n13081), .B(pipeline_rs2_data_bypassed[19]), .S(n9525), 
        .Z(n6313) );
  MUX2_X2 U14600 ( .A(n13082), .B(pipeline_rs2_data_bypassed[20]), .S(n9524), 
        .Z(n6312) );
  MUX2_X2 U14601 ( .A(n13083), .B(pipeline_rs2_data_bypassed[21]), .S(n9523), 
        .Z(n6311) );
  MUX2_X2 U14602 ( .A(n13084), .B(pipeline_rs2_data_bypassed[22]), .S(n9522), 
        .Z(n6310) );
  MUX2_X2 U14603 ( .A(n13085), .B(pipeline_rs2_data_bypassed[23]), .S(n9524), 
        .Z(n6309) );
  MUX2_X2 U14604 ( .A(n13086), .B(pipeline_rs2_data_bypassed[8]), .S(n9525), 
        .Z(n6324) );
  MUX2_X2 U14605 ( .A(n13087), .B(pipeline_rs2_data_bypassed[24]), .S(n9524), 
        .Z(n6308) );
  MUX2_X2 U14606 ( .A(n13088), .B(pipeline_rs2_data_bypassed[9]), .S(n9523), 
        .Z(n6323) );
  MUX2_X2 U14607 ( .A(n13089), .B(pipeline_rs2_data_bypassed[25]), .S(n9523), 
        .Z(n6307) );
  MUX2_X2 U14608 ( .A(n13090), .B(pipeline_rs2_data_bypassed[26]), .S(n9523), 
        .Z(n6306) );
  MUX2_X2 U14609 ( .A(n13091), .B(pipeline_rs2_data_bypassed[27]), .S(n9525), 
        .Z(n6305) );
  MUX2_X2 U14610 ( .A(n13092), .B(pipeline_rs2_data_bypassed[28]), .S(n9522), 
        .Z(n6304) );
  MUX2_X2 U14611 ( .A(n13093), .B(pipeline_rs2_data_bypassed[29]), .S(n9522), 
        .Z(n6303) );
  MUX2_X2 U14612 ( .A(n13094), .B(pipeline_rs2_data_bypassed[30]), .S(n9525), 
        .Z(n6302) );
  MUX2_X2 U14613 ( .A(pipeline_store_data_WB_31_), .B(
        pipeline_rs2_data_bypassed[31]), .S(n9524), .Z(n13136) );
  NAND3_X2 U14614 ( .A1(n9526), .A2(n13099), .A3(n13098), .ZN(n13100) );
  NOR4_X2 U14615 ( .A1(n13100), .A2(n6640), .A3(n9465), .A4(n9527), .ZN(n13121) );
  NOR2_X2 U14616 ( .A1(n13102), .A2(n13101), .ZN(n13107) );
  NAND3_X2 U14617 ( .A1(n13105), .A2(n13104), .A3(n13103), .ZN(n13106) );
  AOI221_X2 U14618 ( .B1(n7181), .B2(n13107), .C1(n7051), .C2(n7081), .A(
        n13106), .ZN(n13120) );
  NOR3_X2 U14619 ( .A1(n13108), .A2(n6697), .A3(n9466), .ZN(n13109) );
  NAND4_X2 U14620 ( .A1(n13112), .A2(n13111), .A3(n13110), .A4(n13109), .ZN(
        n13118) );
  NAND3_X2 U14621 ( .A1(n13115), .A2(n13114), .A3(n13113), .ZN(n13117) );
  NOR4_X2 U14622 ( .A1(n13118), .A2(n13117), .A3(n13116), .A4(n9461), .ZN(
        n13119) );
  NAND3_X2 U14623 ( .A1(n13121), .A2(n13120), .A3(n13119), .ZN(n13122) );
  NAND2_X2 U14624 ( .A1(n8223), .A2(n13122), .ZN(n6370) );
  NOR2_X2 U14625 ( .A1(n10407), .A2(pipeline_inst_DX[29]), .ZN(n13124) );
  NAND2_X2 U14626 ( .A1(pipeline_inst_DX[28]), .A2(n10323), .ZN(n13123) );
  OAI22_X2 U14627 ( .A1(n13124), .A2(n13123), .B1(pipeline_ctrl_N82), .B2(
        n9632), .ZN(pipeline_csr_N79) );
  INV_X4 U14628 ( .A(n13125), .ZN(dmem_hwrite) );
  NOR2_X1 U14629 ( .A1(pipeline_md_N22), .A2(pipeline_md_N21), .ZN(n13133) );
  AOI21_X1 U14630 ( .B1(pipeline_md_N21), .B2(pipeline_md_N22), .A(n13133), 
        .ZN(n13132) );
  NAND2_X1 U14631 ( .A1(n13133), .A2(n13127), .ZN(n13134) );
  OAI21_X1 U14632 ( .B1(n13133), .B2(n13127), .A(n13134), .ZN(pipeline_md_N181) );
  XNOR2_X1 U14633 ( .A(pipeline_md_N24), .B(n13134), .ZN(pipeline_md_N182) );
  NOR2_X1 U14634 ( .A1(pipeline_md_N24), .A2(n13134), .ZN(n13135) );
  XOR2_X1 U14635 ( .A(pipeline_md_N25), .B(n13135), .Z(pipeline_md_N183) );
  NAND2_X2 U14636 ( .A1(n13128), .A2(n6747), .ZN(n13156) );
  NAND3_X2 U14637 ( .A1(n13145), .A2(n13126), .A3(n13127), .ZN(n13152) );
  NOR2_X2 U14638 ( .A1(n13156), .A2(n13152), .ZN(pipeline_md_N315) );
  NAND3_X2 U14639 ( .A1(n13127), .A2(n13126), .A3(pipeline_md_N24), .ZN(n13157) );
  NAND2_X2 U14640 ( .A1(pipeline_md_N22), .A2(n13128), .ZN(n13153) );
  NOR2_X2 U14641 ( .A1(n13157), .A2(n13153), .ZN(pipeline_md_N325) );
  NAND2_X2 U14642 ( .A1(pipeline_md_N22), .A2(pipeline_md_N21), .ZN(n13154) );
  NOR2_X2 U14643 ( .A1(n13157), .A2(n13154), .ZN(pipeline_md_N326) );
  NOR2_X2 U14644 ( .A1(n13127), .A2(n13145), .ZN(n13150) );
  NAND2_X2 U14645 ( .A1(n13150), .A2(n13126), .ZN(n13146) );
  NOR2_X2 U14646 ( .A1(n13156), .A2(n13146), .ZN(pipeline_md_N327) );
  NAND2_X2 U14647 ( .A1(pipeline_md_N21), .A2(n6747), .ZN(n13158) );
  NOR2_X2 U14648 ( .A1(n13158), .A2(n13146), .ZN(pipeline_md_N328) );
  NOR2_X2 U14649 ( .A1(n13153), .A2(n13146), .ZN(pipeline_md_N329) );
  NOR2_X2 U14650 ( .A1(n13154), .A2(n13146), .ZN(pipeline_md_N330) );
  NAND3_X2 U14651 ( .A1(n13127), .A2(n13145), .A3(pipeline_md_N25), .ZN(n13147) );
  NOR2_X2 U14652 ( .A1(n13156), .A2(n13147), .ZN(pipeline_md_N331) );
  NOR2_X2 U14653 ( .A1(n13158), .A2(n13147), .ZN(pipeline_md_N332) );
  NOR2_X2 U14654 ( .A1(n13153), .A2(n13147), .ZN(pipeline_md_N333) );
  NOR2_X2 U14655 ( .A1(n13154), .A2(n13147), .ZN(pipeline_md_N334) );
  NOR2_X2 U14656 ( .A1(n13158), .A2(n13152), .ZN(pipeline_md_N316) );
  NAND3_X2 U14657 ( .A1(pipeline_md_N23), .A2(n13145), .A3(pipeline_md_N25), 
        .ZN(n13148) );
  NOR2_X2 U14658 ( .A1(n13156), .A2(n13148), .ZN(pipeline_md_N335) );
  NOR2_X2 U14659 ( .A1(n13158), .A2(n13148), .ZN(pipeline_md_N336) );
  NOR2_X2 U14660 ( .A1(n13153), .A2(n13148), .ZN(pipeline_md_N337) );
  NOR2_X2 U14661 ( .A1(n13154), .A2(n13148), .ZN(pipeline_md_N338) );
  NAND3_X2 U14662 ( .A1(pipeline_md_N24), .A2(n13127), .A3(pipeline_md_N25), 
        .ZN(n13149) );
  NOR2_X2 U14663 ( .A1(n13156), .A2(n13149), .ZN(pipeline_md_N339) );
  NOR2_X2 U14664 ( .A1(n13158), .A2(n13149), .ZN(pipeline_md_N340) );
  NOR2_X2 U14665 ( .A1(n13153), .A2(n13149), .ZN(pipeline_md_N341) );
  NOR2_X2 U14666 ( .A1(n13154), .A2(n13149), .ZN(pipeline_md_N342) );
  NAND2_X2 U14667 ( .A1(pipeline_md_N25), .A2(n13150), .ZN(n13151) );
  NOR2_X2 U14668 ( .A1(n13156), .A2(n13151), .ZN(pipeline_md_N343) );
  NOR2_X2 U14669 ( .A1(n13158), .A2(n13151), .ZN(pipeline_md_N344) );
  NOR2_X2 U14670 ( .A1(n13153), .A2(n13152), .ZN(pipeline_md_N317) );
  NOR2_X2 U14671 ( .A1(n13153), .A2(n13151), .ZN(pipeline_md_N345) );
  NOR2_X2 U14672 ( .A1(n13154), .A2(n13151), .ZN(pipeline_md_N346) );
  NOR2_X2 U14673 ( .A1(n13154), .A2(n13152), .ZN(pipeline_md_N318) );
  NAND3_X2 U14674 ( .A1(n13145), .A2(n13126), .A3(pipeline_md_N23), .ZN(n13155) );
  NOR2_X2 U14675 ( .A1(n13156), .A2(n13155), .ZN(pipeline_md_N319) );
  NOR2_X2 U14676 ( .A1(n13158), .A2(n13155), .ZN(pipeline_md_N320) );
  NOR2_X2 U14677 ( .A1(n13155), .A2(n13153), .ZN(pipeline_md_N321) );
  NOR2_X2 U14678 ( .A1(n13155), .A2(n13154), .ZN(pipeline_md_N322) );
  NOR2_X2 U14679 ( .A1(n13157), .A2(n13156), .ZN(pipeline_md_N323) );
  NOR2_X2 U14680 ( .A1(n13158), .A2(n13157), .ZN(pipeline_md_N324) );
  INV_X4 U14681 ( .A(n2041), .ZN(n13138) );
  INV_X4 U14682 ( .A(n2042), .ZN(n13139) );
  INV_X4 U14683 ( .A(htif_pcr_req_addr[11]), .ZN(n13140) );
  INV_X4 U14684 ( .A(htif_pcr_req_data[1]), .ZN(n13141) );
  INV_X4 U14685 ( .A(n4229), .ZN(n13143) );
  NAND2_X2 U6097 ( .A1(n10348), .A2(n13130), .ZN(n12827) );
  NAND3_X2 U6098 ( .A1(n7193), .A2(pipeline_regfile_N17), .A3(n9402), .ZN(
        n12615) );
  INV_X4 U6099 ( .A(n9304), .ZN(n9305) );
  NAND3_X2 U6100 ( .A1(pipeline_regfile_N17), .A2(n7166), .A3(n7174), .ZN(
        n11262) );
  INV_X1 U6101 ( .A(n12805), .ZN(n9514) );
  NAND2_X2 U6102 ( .A1(n9398), .A2(n9339), .ZN(n12582) );
  INV_X4 U6103 ( .A(n9322), .ZN(n9323) );
  OAI221_X1 U6104 ( .B1(n416), .B2(n6694), .C1(n475), .C2(n10144), .A(n9779), 
        .ZN(n9780) );
  OAI221_X1 U6105 ( .B1(n426), .B2(n6694), .C1(n480), .C2(n10144), .A(n9754), 
        .ZN(n9755) );
  OAI221_X1 U6106 ( .B1(n422), .B2(n6694), .C1(n478), .C2(n10144), .A(n9782), 
        .ZN(n12944) );
  OAI221_X1 U6107 ( .B1(n454), .B2(n6694), .C1(n494), .C2(n10144), .A(n9752), 
        .ZN(n12870) );
  OAI22_X1 U6108 ( .A1(n12765), .A2(n10159), .B1(n1143), .B2(n12763), .ZN(
        n5709) );
  OAI22_X1 U6109 ( .A1(n12765), .A2(n10160), .B1(n1142), .B2(n12763), .ZN(
        n5708) );
  OAI22_X1 U6110 ( .A1(n12765), .A2(n10161), .B1(n1141), .B2(n12763), .ZN(
        n5707) );
  OAI22_X1 U6111 ( .A1(n12765), .A2(n10162), .B1(n1140), .B2(n12763), .ZN(
        n5706) );
  OAI22_X1 U6112 ( .A1(n1115), .A2(n9504), .B1(n12765), .B2(n10442), .ZN(
        n10443) );
  OAI22_X1 U6113 ( .A1(n13055), .A2(n9504), .B1(n12765), .B2(n10528), .ZN(
        n10529) );
  OAI22_X1 U6114 ( .A1(n1159), .A2(n13105), .B1(n1243), .B2(n11235), .ZN(
        n10900) );
  OAI22_X1 U6115 ( .A1(n1158), .A2(n13105), .B1(n1238), .B2(n11235), .ZN(
        n11117) );
  OAI22_X1 U6116 ( .A1(n13098), .A2(n10998), .B1(n11235), .B2(n10997), .ZN(
        n10999) );
  OAI22_X1 U6117 ( .A1(n11235), .A2(n11234), .B1(n12804), .B2(n11262), .ZN(
        n11236) );
  OAI22_X1 U6118 ( .A1(n1157), .A2(n13105), .B1(n1231), .B2(n11235), .ZN(
        n10627) );
  OAI22_X1 U6119 ( .A1(n13099), .A2(n6866), .B1(n11235), .B2(n10249), .ZN(
        n10250) );
  OAI22_X1 U6120 ( .A1(n13099), .A2(n6845), .B1(n11235), .B2(n10680), .ZN(
        n10681) );
  OAI221_X1 U6121 ( .B1(n6747), .B2(n9521), .C1(n13132), .C2(n13029), .A(
        n13031), .ZN(n6250) );
  OAI22_X1 U6122 ( .A1(n1039), .A2(n9520), .B1(n1040), .B2(n13029), .ZN(n5764)
         );
  OAI22_X1 U6123 ( .A1(n1038), .A2(n9520), .B1(n1039), .B2(n13029), .ZN(n5765)
         );
  OAI22_X1 U6124 ( .A1(n1037), .A2(n9520), .B1(n1038), .B2(n13029), .ZN(n5766)
         );
  OAI22_X1 U6125 ( .A1(n1036), .A2(n9520), .B1(n1037), .B2(n13029), .ZN(n5767)
         );
  OAI22_X1 U6126 ( .A1(n1035), .A2(n9520), .B1(n1036), .B2(n13029), .ZN(n5768)
         );
  OAI22_X1 U6127 ( .A1(n12753), .A2(n10207), .B1(n948), .B2(n6809), .ZN(n5596)
         );
  OAI22_X1 U6128 ( .A1(n12753), .A2(n10208), .B1(n946), .B2(n6809), .ZN(n5597)
         );
  OAI22_X1 U6129 ( .A1(n12753), .A2(n10209), .B1(n944), .B2(n6809), .ZN(n5598)
         );
  OAI22_X1 U6130 ( .A1(n12753), .A2(n10210), .B1(n942), .B2(n6809), .ZN(n5599)
         );
  OAI22_X1 U6131 ( .A1(n12753), .A2(n10211), .B1(n940), .B2(n6809), .ZN(n5600)
         );
  OAI22_X1 U6132 ( .A1(n12753), .A2(n10212), .B1(n938), .B2(n6809), .ZN(n5601)
         );
  OAI22_X1 U6133 ( .A1(n12753), .A2(n10213), .B1(n936), .B2(n6809), .ZN(n5602)
         );
  NAND2_X4 U6134 ( .A1(htif_pcr_req_valid), .A2(htif_pcr_req_ready), .ZN(n2009) );
  INV_X8 U6135 ( .A(n9503), .ZN(n9504) );
endmodule